//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW5AT-LV138PG484AC1/I0
//Device: GW5AT-138
//Device Version: B
//Created Time: Sun May  5 21:58:51 2024

module gowin_data_ram (dout, wre, wad, di, rad, clk);

output [31:0] dout;
input wre;
input [10:0] wad;
input [31:0] di;
input [10:0] rad;
input clk;

wire wad4_inv;
wire wad5_inv;
wire wad6_inv;
wire lut_f_0;
wire wad7_inv;
wire wad8_inv;
wire wad9_inv;
wire wad10_inv;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire lut_f_53;
wire lut_f_54;
wire lut_f_55;
wire lut_f_56;
wire lut_f_57;
wire lut_f_58;
wire lut_f_59;
wire lut_f_60;
wire lut_f_61;
wire lut_f_62;
wire lut_f_63;
wire lut_f_64;
wire lut_f_65;
wire lut_f_66;
wire lut_f_67;
wire lut_f_68;
wire lut_f_69;
wire lut_f_70;
wire lut_f_71;
wire lut_f_72;
wire lut_f_73;
wire lut_f_74;
wire lut_f_75;
wire lut_f_76;
wire lut_f_77;
wire lut_f_78;
wire lut_f_79;
wire lut_f_80;
wire lut_f_81;
wire lut_f_82;
wire lut_f_83;
wire lut_f_84;
wire lut_f_85;
wire lut_f_86;
wire lut_f_87;
wire lut_f_88;
wire lut_f_89;
wire lut_f_90;
wire lut_f_91;
wire lut_f_92;
wire lut_f_93;
wire lut_f_94;
wire lut_f_95;
wire lut_f_96;
wire lut_f_97;
wire lut_f_98;
wire lut_f_99;
wire lut_f_100;
wire lut_f_101;
wire lut_f_102;
wire lut_f_103;
wire lut_f_104;
wire lut_f_105;
wire lut_f_106;
wire lut_f_107;
wire lut_f_108;
wire lut_f_109;
wire lut_f_110;
wire lut_f_111;
wire lut_f_112;
wire lut_f_113;
wire lut_f_114;
wire lut_f_115;
wire lut_f_116;
wire lut_f_117;
wire lut_f_118;
wire lut_f_119;
wire lut_f_120;
wire lut_f_121;
wire lut_f_122;
wire lut_f_123;
wire lut_f_124;
wire lut_f_125;
wire lut_f_126;
wire lut_f_127;
wire lut_f_128;
wire lut_f_129;
wire lut_f_130;
wire lut_f_131;
wire lut_f_132;
wire lut_f_133;
wire lut_f_134;
wire lut_f_135;
wire lut_f_136;
wire lut_f_137;
wire lut_f_138;
wire lut_f_139;
wire lut_f_140;
wire lut_f_141;
wire lut_f_142;
wire lut_f_143;
wire lut_f_144;
wire lut_f_145;
wire lut_f_146;
wire lut_f_147;
wire lut_f_148;
wire lut_f_149;
wire lut_f_150;
wire lut_f_151;
wire lut_f_152;
wire lut_f_153;
wire lut_f_154;
wire lut_f_155;
wire lut_f_156;
wire lut_f_157;
wire lut_f_158;
wire lut_f_159;
wire lut_f_160;
wire lut_f_161;
wire lut_f_162;
wire lut_f_163;
wire lut_f_164;
wire lut_f_165;
wire lut_f_166;
wire lut_f_167;
wire lut_f_168;
wire lut_f_169;
wire lut_f_170;
wire lut_f_171;
wire lut_f_172;
wire lut_f_173;
wire lut_f_174;
wire lut_f_175;
wire lut_f_176;
wire lut_f_177;
wire lut_f_178;
wire lut_f_179;
wire lut_f_180;
wire lut_f_181;
wire lut_f_182;
wire lut_f_183;
wire lut_f_184;
wire lut_f_185;
wire lut_f_186;
wire lut_f_187;
wire lut_f_188;
wire lut_f_189;
wire lut_f_190;
wire lut_f_191;
wire lut_f_192;
wire lut_f_193;
wire lut_f_194;
wire lut_f_195;
wire lut_f_196;
wire lut_f_197;
wire lut_f_198;
wire lut_f_199;
wire lut_f_200;
wire lut_f_201;
wire lut_f_202;
wire lut_f_203;
wire lut_f_204;
wire lut_f_205;
wire lut_f_206;
wire lut_f_207;
wire lut_f_208;
wire lut_f_209;
wire lut_f_210;
wire lut_f_211;
wire lut_f_212;
wire lut_f_213;
wire lut_f_214;
wire lut_f_215;
wire lut_f_216;
wire lut_f_217;
wire lut_f_218;
wire lut_f_219;
wire lut_f_220;
wire lut_f_221;
wire lut_f_222;
wire lut_f_223;
wire lut_f_224;
wire lut_f_225;
wire lut_f_226;
wire lut_f_227;
wire lut_f_228;
wire lut_f_229;
wire lut_f_230;
wire lut_f_231;
wire lut_f_232;
wire lut_f_233;
wire lut_f_234;
wire lut_f_235;
wire lut_f_236;
wire lut_f_237;
wire lut_f_238;
wire lut_f_239;
wire lut_f_240;
wire lut_f_241;
wire lut_f_242;
wire lut_f_243;
wire lut_f_244;
wire lut_f_245;
wire lut_f_246;
wire lut_f_247;
wire lut_f_248;
wire lut_f_249;
wire lut_f_250;
wire lut_f_251;
wire lut_f_252;
wire lut_f_253;
wire lut_f_254;
wire lut_f_255;
wire lut_f_256;
wire lut_f_257;
wire lut_f_258;
wire lut_f_259;
wire lut_f_260;
wire lut_f_261;
wire lut_f_262;
wire lut_f_263;
wire lut_f_264;
wire lut_f_265;
wire lut_f_266;
wire lut_f_267;
wire lut_f_268;
wire lut_f_269;
wire lut_f_270;
wire lut_f_271;
wire lut_f_272;
wire lut_f_273;
wire lut_f_274;
wire lut_f_275;
wire lut_f_276;
wire lut_f_277;
wire lut_f_278;
wire lut_f_279;
wire lut_f_280;
wire lut_f_281;
wire lut_f_282;
wire lut_f_283;
wire lut_f_284;
wire lut_f_285;
wire lut_f_286;
wire lut_f_287;
wire lut_f_288;
wire lut_f_289;
wire lut_f_290;
wire lut_f_291;
wire lut_f_292;
wire lut_f_293;
wire lut_f_294;
wire lut_f_295;
wire lut_f_296;
wire lut_f_297;
wire lut_f_298;
wire lut_f_299;
wire lut_f_300;
wire lut_f_301;
wire lut_f_302;
wire lut_f_303;
wire lut_f_304;
wire lut_f_305;
wire lut_f_306;
wire lut_f_307;
wire lut_f_308;
wire lut_f_309;
wire lut_f_310;
wire lut_f_311;
wire lut_f_312;
wire lut_f_313;
wire lut_f_314;
wire lut_f_315;
wire lut_f_316;
wire lut_f_317;
wire lut_f_318;
wire lut_f_319;
wire lut_f_320;
wire lut_f_321;
wire lut_f_322;
wire lut_f_323;
wire lut_f_324;
wire lut_f_325;
wire lut_f_326;
wire lut_f_327;
wire lut_f_328;
wire lut_f_329;
wire lut_f_330;
wire lut_f_331;
wire lut_f_332;
wire lut_f_333;
wire lut_f_334;
wire lut_f_335;
wire lut_f_336;
wire lut_f_337;
wire lut_f_338;
wire lut_f_339;
wire lut_f_340;
wire lut_f_341;
wire lut_f_342;
wire lut_f_343;
wire lut_f_344;
wire lut_f_345;
wire lut_f_346;
wire lut_f_347;
wire lut_f_348;
wire lut_f_349;
wire lut_f_350;
wire lut_f_351;
wire lut_f_352;
wire lut_f_353;
wire lut_f_354;
wire lut_f_355;
wire lut_f_356;
wire lut_f_357;
wire lut_f_358;
wire lut_f_359;
wire lut_f_360;
wire lut_f_361;
wire lut_f_362;
wire lut_f_363;
wire lut_f_364;
wire lut_f_365;
wire lut_f_366;
wire lut_f_367;
wire lut_f_368;
wire lut_f_369;
wire lut_f_370;
wire lut_f_371;
wire lut_f_372;
wire lut_f_373;
wire lut_f_374;
wire lut_f_375;
wire lut_f_376;
wire lut_f_377;
wire lut_f_378;
wire lut_f_379;
wire lut_f_380;
wire lut_f_381;
wire lut_f_382;
wire lut_f_383;
wire [3:0] ram16sdp_inst_0_dout;
wire [7:4] ram16sdp_inst_1_dout;
wire [11:8] ram16sdp_inst_2_dout;
wire [15:12] ram16sdp_inst_3_dout;
wire [19:16] ram16sdp_inst_4_dout;
wire [23:20] ram16sdp_inst_5_dout;
wire [27:24] ram16sdp_inst_6_dout;
wire [31:28] ram16sdp_inst_7_dout;
wire [3:0] ram16sdp_inst_8_dout;
wire [7:4] ram16sdp_inst_9_dout;
wire [11:8] ram16sdp_inst_10_dout;
wire [15:12] ram16sdp_inst_11_dout;
wire [19:16] ram16sdp_inst_12_dout;
wire [23:20] ram16sdp_inst_13_dout;
wire [27:24] ram16sdp_inst_14_dout;
wire [31:28] ram16sdp_inst_15_dout;
wire [3:0] ram16sdp_inst_16_dout;
wire [7:4] ram16sdp_inst_17_dout;
wire [11:8] ram16sdp_inst_18_dout;
wire [15:12] ram16sdp_inst_19_dout;
wire [19:16] ram16sdp_inst_20_dout;
wire [23:20] ram16sdp_inst_21_dout;
wire [27:24] ram16sdp_inst_22_dout;
wire [31:28] ram16sdp_inst_23_dout;
wire [3:0] ram16sdp_inst_24_dout;
wire [7:4] ram16sdp_inst_25_dout;
wire [11:8] ram16sdp_inst_26_dout;
wire [15:12] ram16sdp_inst_27_dout;
wire [19:16] ram16sdp_inst_28_dout;
wire [23:20] ram16sdp_inst_29_dout;
wire [27:24] ram16sdp_inst_30_dout;
wire [31:28] ram16sdp_inst_31_dout;
wire [3:0] ram16sdp_inst_32_dout;
wire [7:4] ram16sdp_inst_33_dout;
wire [11:8] ram16sdp_inst_34_dout;
wire [15:12] ram16sdp_inst_35_dout;
wire [19:16] ram16sdp_inst_36_dout;
wire [23:20] ram16sdp_inst_37_dout;
wire [27:24] ram16sdp_inst_38_dout;
wire [31:28] ram16sdp_inst_39_dout;
wire [3:0] ram16sdp_inst_40_dout;
wire [7:4] ram16sdp_inst_41_dout;
wire [11:8] ram16sdp_inst_42_dout;
wire [15:12] ram16sdp_inst_43_dout;
wire [19:16] ram16sdp_inst_44_dout;
wire [23:20] ram16sdp_inst_45_dout;
wire [27:24] ram16sdp_inst_46_dout;
wire [31:28] ram16sdp_inst_47_dout;
wire [3:0] ram16sdp_inst_48_dout;
wire [7:4] ram16sdp_inst_49_dout;
wire [11:8] ram16sdp_inst_50_dout;
wire [15:12] ram16sdp_inst_51_dout;
wire [19:16] ram16sdp_inst_52_dout;
wire [23:20] ram16sdp_inst_53_dout;
wire [27:24] ram16sdp_inst_54_dout;
wire [31:28] ram16sdp_inst_55_dout;
wire [3:0] ram16sdp_inst_56_dout;
wire [7:4] ram16sdp_inst_57_dout;
wire [11:8] ram16sdp_inst_58_dout;
wire [15:12] ram16sdp_inst_59_dout;
wire [19:16] ram16sdp_inst_60_dout;
wire [23:20] ram16sdp_inst_61_dout;
wire [27:24] ram16sdp_inst_62_dout;
wire [31:28] ram16sdp_inst_63_dout;
wire [3:0] ram16sdp_inst_64_dout;
wire [7:4] ram16sdp_inst_65_dout;
wire [11:8] ram16sdp_inst_66_dout;
wire [15:12] ram16sdp_inst_67_dout;
wire [19:16] ram16sdp_inst_68_dout;
wire [23:20] ram16sdp_inst_69_dout;
wire [27:24] ram16sdp_inst_70_dout;
wire [31:28] ram16sdp_inst_71_dout;
wire [3:0] ram16sdp_inst_72_dout;
wire [7:4] ram16sdp_inst_73_dout;
wire [11:8] ram16sdp_inst_74_dout;
wire [15:12] ram16sdp_inst_75_dout;
wire [19:16] ram16sdp_inst_76_dout;
wire [23:20] ram16sdp_inst_77_dout;
wire [27:24] ram16sdp_inst_78_dout;
wire [31:28] ram16sdp_inst_79_dout;
wire [3:0] ram16sdp_inst_80_dout;
wire [7:4] ram16sdp_inst_81_dout;
wire [11:8] ram16sdp_inst_82_dout;
wire [15:12] ram16sdp_inst_83_dout;
wire [19:16] ram16sdp_inst_84_dout;
wire [23:20] ram16sdp_inst_85_dout;
wire [27:24] ram16sdp_inst_86_dout;
wire [31:28] ram16sdp_inst_87_dout;
wire [3:0] ram16sdp_inst_88_dout;
wire [7:4] ram16sdp_inst_89_dout;
wire [11:8] ram16sdp_inst_90_dout;
wire [15:12] ram16sdp_inst_91_dout;
wire [19:16] ram16sdp_inst_92_dout;
wire [23:20] ram16sdp_inst_93_dout;
wire [27:24] ram16sdp_inst_94_dout;
wire [31:28] ram16sdp_inst_95_dout;
wire [3:0] ram16sdp_inst_96_dout;
wire [7:4] ram16sdp_inst_97_dout;
wire [11:8] ram16sdp_inst_98_dout;
wire [15:12] ram16sdp_inst_99_dout;
wire [19:16] ram16sdp_inst_100_dout;
wire [23:20] ram16sdp_inst_101_dout;
wire [27:24] ram16sdp_inst_102_dout;
wire [31:28] ram16sdp_inst_103_dout;
wire [3:0] ram16sdp_inst_104_dout;
wire [7:4] ram16sdp_inst_105_dout;
wire [11:8] ram16sdp_inst_106_dout;
wire [15:12] ram16sdp_inst_107_dout;
wire [19:16] ram16sdp_inst_108_dout;
wire [23:20] ram16sdp_inst_109_dout;
wire [27:24] ram16sdp_inst_110_dout;
wire [31:28] ram16sdp_inst_111_dout;
wire [3:0] ram16sdp_inst_112_dout;
wire [7:4] ram16sdp_inst_113_dout;
wire [11:8] ram16sdp_inst_114_dout;
wire [15:12] ram16sdp_inst_115_dout;
wire [19:16] ram16sdp_inst_116_dout;
wire [23:20] ram16sdp_inst_117_dout;
wire [27:24] ram16sdp_inst_118_dout;
wire [31:28] ram16sdp_inst_119_dout;
wire [3:0] ram16sdp_inst_120_dout;
wire [7:4] ram16sdp_inst_121_dout;
wire [11:8] ram16sdp_inst_122_dout;
wire [15:12] ram16sdp_inst_123_dout;
wire [19:16] ram16sdp_inst_124_dout;
wire [23:20] ram16sdp_inst_125_dout;
wire [27:24] ram16sdp_inst_126_dout;
wire [31:28] ram16sdp_inst_127_dout;
wire [3:0] ram16sdp_inst_128_dout;
wire [7:4] ram16sdp_inst_129_dout;
wire [11:8] ram16sdp_inst_130_dout;
wire [15:12] ram16sdp_inst_131_dout;
wire [19:16] ram16sdp_inst_132_dout;
wire [23:20] ram16sdp_inst_133_dout;
wire [27:24] ram16sdp_inst_134_dout;
wire [31:28] ram16sdp_inst_135_dout;
wire [3:0] ram16sdp_inst_136_dout;
wire [7:4] ram16sdp_inst_137_dout;
wire [11:8] ram16sdp_inst_138_dout;
wire [15:12] ram16sdp_inst_139_dout;
wire [19:16] ram16sdp_inst_140_dout;
wire [23:20] ram16sdp_inst_141_dout;
wire [27:24] ram16sdp_inst_142_dout;
wire [31:28] ram16sdp_inst_143_dout;
wire [3:0] ram16sdp_inst_144_dout;
wire [7:4] ram16sdp_inst_145_dout;
wire [11:8] ram16sdp_inst_146_dout;
wire [15:12] ram16sdp_inst_147_dout;
wire [19:16] ram16sdp_inst_148_dout;
wire [23:20] ram16sdp_inst_149_dout;
wire [27:24] ram16sdp_inst_150_dout;
wire [31:28] ram16sdp_inst_151_dout;
wire [3:0] ram16sdp_inst_152_dout;
wire [7:4] ram16sdp_inst_153_dout;
wire [11:8] ram16sdp_inst_154_dout;
wire [15:12] ram16sdp_inst_155_dout;
wire [19:16] ram16sdp_inst_156_dout;
wire [23:20] ram16sdp_inst_157_dout;
wire [27:24] ram16sdp_inst_158_dout;
wire [31:28] ram16sdp_inst_159_dout;
wire [3:0] ram16sdp_inst_160_dout;
wire [7:4] ram16sdp_inst_161_dout;
wire [11:8] ram16sdp_inst_162_dout;
wire [15:12] ram16sdp_inst_163_dout;
wire [19:16] ram16sdp_inst_164_dout;
wire [23:20] ram16sdp_inst_165_dout;
wire [27:24] ram16sdp_inst_166_dout;
wire [31:28] ram16sdp_inst_167_dout;
wire [3:0] ram16sdp_inst_168_dout;
wire [7:4] ram16sdp_inst_169_dout;
wire [11:8] ram16sdp_inst_170_dout;
wire [15:12] ram16sdp_inst_171_dout;
wire [19:16] ram16sdp_inst_172_dout;
wire [23:20] ram16sdp_inst_173_dout;
wire [27:24] ram16sdp_inst_174_dout;
wire [31:28] ram16sdp_inst_175_dout;
wire [3:0] ram16sdp_inst_176_dout;
wire [7:4] ram16sdp_inst_177_dout;
wire [11:8] ram16sdp_inst_178_dout;
wire [15:12] ram16sdp_inst_179_dout;
wire [19:16] ram16sdp_inst_180_dout;
wire [23:20] ram16sdp_inst_181_dout;
wire [27:24] ram16sdp_inst_182_dout;
wire [31:28] ram16sdp_inst_183_dout;
wire [3:0] ram16sdp_inst_184_dout;
wire [7:4] ram16sdp_inst_185_dout;
wire [11:8] ram16sdp_inst_186_dout;
wire [15:12] ram16sdp_inst_187_dout;
wire [19:16] ram16sdp_inst_188_dout;
wire [23:20] ram16sdp_inst_189_dout;
wire [27:24] ram16sdp_inst_190_dout;
wire [31:28] ram16sdp_inst_191_dout;
wire [3:0] ram16sdp_inst_192_dout;
wire [7:4] ram16sdp_inst_193_dout;
wire [11:8] ram16sdp_inst_194_dout;
wire [15:12] ram16sdp_inst_195_dout;
wire [19:16] ram16sdp_inst_196_dout;
wire [23:20] ram16sdp_inst_197_dout;
wire [27:24] ram16sdp_inst_198_dout;
wire [31:28] ram16sdp_inst_199_dout;
wire [3:0] ram16sdp_inst_200_dout;
wire [7:4] ram16sdp_inst_201_dout;
wire [11:8] ram16sdp_inst_202_dout;
wire [15:12] ram16sdp_inst_203_dout;
wire [19:16] ram16sdp_inst_204_dout;
wire [23:20] ram16sdp_inst_205_dout;
wire [27:24] ram16sdp_inst_206_dout;
wire [31:28] ram16sdp_inst_207_dout;
wire [3:0] ram16sdp_inst_208_dout;
wire [7:4] ram16sdp_inst_209_dout;
wire [11:8] ram16sdp_inst_210_dout;
wire [15:12] ram16sdp_inst_211_dout;
wire [19:16] ram16sdp_inst_212_dout;
wire [23:20] ram16sdp_inst_213_dout;
wire [27:24] ram16sdp_inst_214_dout;
wire [31:28] ram16sdp_inst_215_dout;
wire [3:0] ram16sdp_inst_216_dout;
wire [7:4] ram16sdp_inst_217_dout;
wire [11:8] ram16sdp_inst_218_dout;
wire [15:12] ram16sdp_inst_219_dout;
wire [19:16] ram16sdp_inst_220_dout;
wire [23:20] ram16sdp_inst_221_dout;
wire [27:24] ram16sdp_inst_222_dout;
wire [31:28] ram16sdp_inst_223_dout;
wire [3:0] ram16sdp_inst_224_dout;
wire [7:4] ram16sdp_inst_225_dout;
wire [11:8] ram16sdp_inst_226_dout;
wire [15:12] ram16sdp_inst_227_dout;
wire [19:16] ram16sdp_inst_228_dout;
wire [23:20] ram16sdp_inst_229_dout;
wire [27:24] ram16sdp_inst_230_dout;
wire [31:28] ram16sdp_inst_231_dout;
wire [3:0] ram16sdp_inst_232_dout;
wire [7:4] ram16sdp_inst_233_dout;
wire [11:8] ram16sdp_inst_234_dout;
wire [15:12] ram16sdp_inst_235_dout;
wire [19:16] ram16sdp_inst_236_dout;
wire [23:20] ram16sdp_inst_237_dout;
wire [27:24] ram16sdp_inst_238_dout;
wire [31:28] ram16sdp_inst_239_dout;
wire [3:0] ram16sdp_inst_240_dout;
wire [7:4] ram16sdp_inst_241_dout;
wire [11:8] ram16sdp_inst_242_dout;
wire [15:12] ram16sdp_inst_243_dout;
wire [19:16] ram16sdp_inst_244_dout;
wire [23:20] ram16sdp_inst_245_dout;
wire [27:24] ram16sdp_inst_246_dout;
wire [31:28] ram16sdp_inst_247_dout;
wire [3:0] ram16sdp_inst_248_dout;
wire [7:4] ram16sdp_inst_249_dout;
wire [11:8] ram16sdp_inst_250_dout;
wire [15:12] ram16sdp_inst_251_dout;
wire [19:16] ram16sdp_inst_252_dout;
wire [23:20] ram16sdp_inst_253_dout;
wire [27:24] ram16sdp_inst_254_dout;
wire [31:28] ram16sdp_inst_255_dout;
wire [3:0] ram16sdp_inst_256_dout;
wire [7:4] ram16sdp_inst_257_dout;
wire [11:8] ram16sdp_inst_258_dout;
wire [15:12] ram16sdp_inst_259_dout;
wire [19:16] ram16sdp_inst_260_dout;
wire [23:20] ram16sdp_inst_261_dout;
wire [27:24] ram16sdp_inst_262_dout;
wire [31:28] ram16sdp_inst_263_dout;
wire [3:0] ram16sdp_inst_264_dout;
wire [7:4] ram16sdp_inst_265_dout;
wire [11:8] ram16sdp_inst_266_dout;
wire [15:12] ram16sdp_inst_267_dout;
wire [19:16] ram16sdp_inst_268_dout;
wire [23:20] ram16sdp_inst_269_dout;
wire [27:24] ram16sdp_inst_270_dout;
wire [31:28] ram16sdp_inst_271_dout;
wire [3:0] ram16sdp_inst_272_dout;
wire [7:4] ram16sdp_inst_273_dout;
wire [11:8] ram16sdp_inst_274_dout;
wire [15:12] ram16sdp_inst_275_dout;
wire [19:16] ram16sdp_inst_276_dout;
wire [23:20] ram16sdp_inst_277_dout;
wire [27:24] ram16sdp_inst_278_dout;
wire [31:28] ram16sdp_inst_279_dout;
wire [3:0] ram16sdp_inst_280_dout;
wire [7:4] ram16sdp_inst_281_dout;
wire [11:8] ram16sdp_inst_282_dout;
wire [15:12] ram16sdp_inst_283_dout;
wire [19:16] ram16sdp_inst_284_dout;
wire [23:20] ram16sdp_inst_285_dout;
wire [27:24] ram16sdp_inst_286_dout;
wire [31:28] ram16sdp_inst_287_dout;
wire [3:0] ram16sdp_inst_288_dout;
wire [7:4] ram16sdp_inst_289_dout;
wire [11:8] ram16sdp_inst_290_dout;
wire [15:12] ram16sdp_inst_291_dout;
wire [19:16] ram16sdp_inst_292_dout;
wire [23:20] ram16sdp_inst_293_dout;
wire [27:24] ram16sdp_inst_294_dout;
wire [31:28] ram16sdp_inst_295_dout;
wire [3:0] ram16sdp_inst_296_dout;
wire [7:4] ram16sdp_inst_297_dout;
wire [11:8] ram16sdp_inst_298_dout;
wire [15:12] ram16sdp_inst_299_dout;
wire [19:16] ram16sdp_inst_300_dout;
wire [23:20] ram16sdp_inst_301_dout;
wire [27:24] ram16sdp_inst_302_dout;
wire [31:28] ram16sdp_inst_303_dout;
wire [3:0] ram16sdp_inst_304_dout;
wire [7:4] ram16sdp_inst_305_dout;
wire [11:8] ram16sdp_inst_306_dout;
wire [15:12] ram16sdp_inst_307_dout;
wire [19:16] ram16sdp_inst_308_dout;
wire [23:20] ram16sdp_inst_309_dout;
wire [27:24] ram16sdp_inst_310_dout;
wire [31:28] ram16sdp_inst_311_dout;
wire [3:0] ram16sdp_inst_312_dout;
wire [7:4] ram16sdp_inst_313_dout;
wire [11:8] ram16sdp_inst_314_dout;
wire [15:12] ram16sdp_inst_315_dout;
wire [19:16] ram16sdp_inst_316_dout;
wire [23:20] ram16sdp_inst_317_dout;
wire [27:24] ram16sdp_inst_318_dout;
wire [31:28] ram16sdp_inst_319_dout;
wire [3:0] ram16sdp_inst_320_dout;
wire [7:4] ram16sdp_inst_321_dout;
wire [11:8] ram16sdp_inst_322_dout;
wire [15:12] ram16sdp_inst_323_dout;
wire [19:16] ram16sdp_inst_324_dout;
wire [23:20] ram16sdp_inst_325_dout;
wire [27:24] ram16sdp_inst_326_dout;
wire [31:28] ram16sdp_inst_327_dout;
wire [3:0] ram16sdp_inst_328_dout;
wire [7:4] ram16sdp_inst_329_dout;
wire [11:8] ram16sdp_inst_330_dout;
wire [15:12] ram16sdp_inst_331_dout;
wire [19:16] ram16sdp_inst_332_dout;
wire [23:20] ram16sdp_inst_333_dout;
wire [27:24] ram16sdp_inst_334_dout;
wire [31:28] ram16sdp_inst_335_dout;
wire [3:0] ram16sdp_inst_336_dout;
wire [7:4] ram16sdp_inst_337_dout;
wire [11:8] ram16sdp_inst_338_dout;
wire [15:12] ram16sdp_inst_339_dout;
wire [19:16] ram16sdp_inst_340_dout;
wire [23:20] ram16sdp_inst_341_dout;
wire [27:24] ram16sdp_inst_342_dout;
wire [31:28] ram16sdp_inst_343_dout;
wire [3:0] ram16sdp_inst_344_dout;
wire [7:4] ram16sdp_inst_345_dout;
wire [11:8] ram16sdp_inst_346_dout;
wire [15:12] ram16sdp_inst_347_dout;
wire [19:16] ram16sdp_inst_348_dout;
wire [23:20] ram16sdp_inst_349_dout;
wire [27:24] ram16sdp_inst_350_dout;
wire [31:28] ram16sdp_inst_351_dout;
wire [3:0] ram16sdp_inst_352_dout;
wire [7:4] ram16sdp_inst_353_dout;
wire [11:8] ram16sdp_inst_354_dout;
wire [15:12] ram16sdp_inst_355_dout;
wire [19:16] ram16sdp_inst_356_dout;
wire [23:20] ram16sdp_inst_357_dout;
wire [27:24] ram16sdp_inst_358_dout;
wire [31:28] ram16sdp_inst_359_dout;
wire [3:0] ram16sdp_inst_360_dout;
wire [7:4] ram16sdp_inst_361_dout;
wire [11:8] ram16sdp_inst_362_dout;
wire [15:12] ram16sdp_inst_363_dout;
wire [19:16] ram16sdp_inst_364_dout;
wire [23:20] ram16sdp_inst_365_dout;
wire [27:24] ram16sdp_inst_366_dout;
wire [31:28] ram16sdp_inst_367_dout;
wire [3:0] ram16sdp_inst_368_dout;
wire [7:4] ram16sdp_inst_369_dout;
wire [11:8] ram16sdp_inst_370_dout;
wire [15:12] ram16sdp_inst_371_dout;
wire [19:16] ram16sdp_inst_372_dout;
wire [23:20] ram16sdp_inst_373_dout;
wire [27:24] ram16sdp_inst_374_dout;
wire [31:28] ram16sdp_inst_375_dout;
wire [3:0] ram16sdp_inst_376_dout;
wire [7:4] ram16sdp_inst_377_dout;
wire [11:8] ram16sdp_inst_378_dout;
wire [15:12] ram16sdp_inst_379_dout;
wire [19:16] ram16sdp_inst_380_dout;
wire [23:20] ram16sdp_inst_381_dout;
wire [27:24] ram16sdp_inst_382_dout;
wire [31:28] ram16sdp_inst_383_dout;
wire [3:0] ram16sdp_inst_384_dout;
wire [7:4] ram16sdp_inst_385_dout;
wire [11:8] ram16sdp_inst_386_dout;
wire [15:12] ram16sdp_inst_387_dout;
wire [19:16] ram16sdp_inst_388_dout;
wire [23:20] ram16sdp_inst_389_dout;
wire [27:24] ram16sdp_inst_390_dout;
wire [31:28] ram16sdp_inst_391_dout;
wire [3:0] ram16sdp_inst_392_dout;
wire [7:4] ram16sdp_inst_393_dout;
wire [11:8] ram16sdp_inst_394_dout;
wire [15:12] ram16sdp_inst_395_dout;
wire [19:16] ram16sdp_inst_396_dout;
wire [23:20] ram16sdp_inst_397_dout;
wire [27:24] ram16sdp_inst_398_dout;
wire [31:28] ram16sdp_inst_399_dout;
wire [3:0] ram16sdp_inst_400_dout;
wire [7:4] ram16sdp_inst_401_dout;
wire [11:8] ram16sdp_inst_402_dout;
wire [15:12] ram16sdp_inst_403_dout;
wire [19:16] ram16sdp_inst_404_dout;
wire [23:20] ram16sdp_inst_405_dout;
wire [27:24] ram16sdp_inst_406_dout;
wire [31:28] ram16sdp_inst_407_dout;
wire [3:0] ram16sdp_inst_408_dout;
wire [7:4] ram16sdp_inst_409_dout;
wire [11:8] ram16sdp_inst_410_dout;
wire [15:12] ram16sdp_inst_411_dout;
wire [19:16] ram16sdp_inst_412_dout;
wire [23:20] ram16sdp_inst_413_dout;
wire [27:24] ram16sdp_inst_414_dout;
wire [31:28] ram16sdp_inst_415_dout;
wire [3:0] ram16sdp_inst_416_dout;
wire [7:4] ram16sdp_inst_417_dout;
wire [11:8] ram16sdp_inst_418_dout;
wire [15:12] ram16sdp_inst_419_dout;
wire [19:16] ram16sdp_inst_420_dout;
wire [23:20] ram16sdp_inst_421_dout;
wire [27:24] ram16sdp_inst_422_dout;
wire [31:28] ram16sdp_inst_423_dout;
wire [3:0] ram16sdp_inst_424_dout;
wire [7:4] ram16sdp_inst_425_dout;
wire [11:8] ram16sdp_inst_426_dout;
wire [15:12] ram16sdp_inst_427_dout;
wire [19:16] ram16sdp_inst_428_dout;
wire [23:20] ram16sdp_inst_429_dout;
wire [27:24] ram16sdp_inst_430_dout;
wire [31:28] ram16sdp_inst_431_dout;
wire [3:0] ram16sdp_inst_432_dout;
wire [7:4] ram16sdp_inst_433_dout;
wire [11:8] ram16sdp_inst_434_dout;
wire [15:12] ram16sdp_inst_435_dout;
wire [19:16] ram16sdp_inst_436_dout;
wire [23:20] ram16sdp_inst_437_dout;
wire [27:24] ram16sdp_inst_438_dout;
wire [31:28] ram16sdp_inst_439_dout;
wire [3:0] ram16sdp_inst_440_dout;
wire [7:4] ram16sdp_inst_441_dout;
wire [11:8] ram16sdp_inst_442_dout;
wire [15:12] ram16sdp_inst_443_dout;
wire [19:16] ram16sdp_inst_444_dout;
wire [23:20] ram16sdp_inst_445_dout;
wire [27:24] ram16sdp_inst_446_dout;
wire [31:28] ram16sdp_inst_447_dout;
wire [3:0] ram16sdp_inst_448_dout;
wire [7:4] ram16sdp_inst_449_dout;
wire [11:8] ram16sdp_inst_450_dout;
wire [15:12] ram16sdp_inst_451_dout;
wire [19:16] ram16sdp_inst_452_dout;
wire [23:20] ram16sdp_inst_453_dout;
wire [27:24] ram16sdp_inst_454_dout;
wire [31:28] ram16sdp_inst_455_dout;
wire [3:0] ram16sdp_inst_456_dout;
wire [7:4] ram16sdp_inst_457_dout;
wire [11:8] ram16sdp_inst_458_dout;
wire [15:12] ram16sdp_inst_459_dout;
wire [19:16] ram16sdp_inst_460_dout;
wire [23:20] ram16sdp_inst_461_dout;
wire [27:24] ram16sdp_inst_462_dout;
wire [31:28] ram16sdp_inst_463_dout;
wire [3:0] ram16sdp_inst_464_dout;
wire [7:4] ram16sdp_inst_465_dout;
wire [11:8] ram16sdp_inst_466_dout;
wire [15:12] ram16sdp_inst_467_dout;
wire [19:16] ram16sdp_inst_468_dout;
wire [23:20] ram16sdp_inst_469_dout;
wire [27:24] ram16sdp_inst_470_dout;
wire [31:28] ram16sdp_inst_471_dout;
wire [3:0] ram16sdp_inst_472_dout;
wire [7:4] ram16sdp_inst_473_dout;
wire [11:8] ram16sdp_inst_474_dout;
wire [15:12] ram16sdp_inst_475_dout;
wire [19:16] ram16sdp_inst_476_dout;
wire [23:20] ram16sdp_inst_477_dout;
wire [27:24] ram16sdp_inst_478_dout;
wire [31:28] ram16sdp_inst_479_dout;
wire [3:0] ram16sdp_inst_480_dout;
wire [7:4] ram16sdp_inst_481_dout;
wire [11:8] ram16sdp_inst_482_dout;
wire [15:12] ram16sdp_inst_483_dout;
wire [19:16] ram16sdp_inst_484_dout;
wire [23:20] ram16sdp_inst_485_dout;
wire [27:24] ram16sdp_inst_486_dout;
wire [31:28] ram16sdp_inst_487_dout;
wire [3:0] ram16sdp_inst_488_dout;
wire [7:4] ram16sdp_inst_489_dout;
wire [11:8] ram16sdp_inst_490_dout;
wire [15:12] ram16sdp_inst_491_dout;
wire [19:16] ram16sdp_inst_492_dout;
wire [23:20] ram16sdp_inst_493_dout;
wire [27:24] ram16sdp_inst_494_dout;
wire [31:28] ram16sdp_inst_495_dout;
wire [3:0] ram16sdp_inst_496_dout;
wire [7:4] ram16sdp_inst_497_dout;
wire [11:8] ram16sdp_inst_498_dout;
wire [15:12] ram16sdp_inst_499_dout;
wire [19:16] ram16sdp_inst_500_dout;
wire [23:20] ram16sdp_inst_501_dout;
wire [27:24] ram16sdp_inst_502_dout;
wire [31:28] ram16sdp_inst_503_dout;
wire [3:0] ram16sdp_inst_504_dout;
wire [7:4] ram16sdp_inst_505_dout;
wire [11:8] ram16sdp_inst_506_dout;
wire [15:12] ram16sdp_inst_507_dout;
wire [19:16] ram16sdp_inst_508_dout;
wire [23:20] ram16sdp_inst_509_dout;
wire [27:24] ram16sdp_inst_510_dout;
wire [31:28] ram16sdp_inst_511_dout;
wire [3:0] ram16sdp_inst_512_dout;
wire [7:4] ram16sdp_inst_513_dout;
wire [11:8] ram16sdp_inst_514_dout;
wire [15:12] ram16sdp_inst_515_dout;
wire [19:16] ram16sdp_inst_516_dout;
wire [23:20] ram16sdp_inst_517_dout;
wire [27:24] ram16sdp_inst_518_dout;
wire [31:28] ram16sdp_inst_519_dout;
wire [3:0] ram16sdp_inst_520_dout;
wire [7:4] ram16sdp_inst_521_dout;
wire [11:8] ram16sdp_inst_522_dout;
wire [15:12] ram16sdp_inst_523_dout;
wire [19:16] ram16sdp_inst_524_dout;
wire [23:20] ram16sdp_inst_525_dout;
wire [27:24] ram16sdp_inst_526_dout;
wire [31:28] ram16sdp_inst_527_dout;
wire [3:0] ram16sdp_inst_528_dout;
wire [7:4] ram16sdp_inst_529_dout;
wire [11:8] ram16sdp_inst_530_dout;
wire [15:12] ram16sdp_inst_531_dout;
wire [19:16] ram16sdp_inst_532_dout;
wire [23:20] ram16sdp_inst_533_dout;
wire [27:24] ram16sdp_inst_534_dout;
wire [31:28] ram16sdp_inst_535_dout;
wire [3:0] ram16sdp_inst_536_dout;
wire [7:4] ram16sdp_inst_537_dout;
wire [11:8] ram16sdp_inst_538_dout;
wire [15:12] ram16sdp_inst_539_dout;
wire [19:16] ram16sdp_inst_540_dout;
wire [23:20] ram16sdp_inst_541_dout;
wire [27:24] ram16sdp_inst_542_dout;
wire [31:28] ram16sdp_inst_543_dout;
wire [3:0] ram16sdp_inst_544_dout;
wire [7:4] ram16sdp_inst_545_dout;
wire [11:8] ram16sdp_inst_546_dout;
wire [15:12] ram16sdp_inst_547_dout;
wire [19:16] ram16sdp_inst_548_dout;
wire [23:20] ram16sdp_inst_549_dout;
wire [27:24] ram16sdp_inst_550_dout;
wire [31:28] ram16sdp_inst_551_dout;
wire [3:0] ram16sdp_inst_552_dout;
wire [7:4] ram16sdp_inst_553_dout;
wire [11:8] ram16sdp_inst_554_dout;
wire [15:12] ram16sdp_inst_555_dout;
wire [19:16] ram16sdp_inst_556_dout;
wire [23:20] ram16sdp_inst_557_dout;
wire [27:24] ram16sdp_inst_558_dout;
wire [31:28] ram16sdp_inst_559_dout;
wire [3:0] ram16sdp_inst_560_dout;
wire [7:4] ram16sdp_inst_561_dout;
wire [11:8] ram16sdp_inst_562_dout;
wire [15:12] ram16sdp_inst_563_dout;
wire [19:16] ram16sdp_inst_564_dout;
wire [23:20] ram16sdp_inst_565_dout;
wire [27:24] ram16sdp_inst_566_dout;
wire [31:28] ram16sdp_inst_567_dout;
wire [3:0] ram16sdp_inst_568_dout;
wire [7:4] ram16sdp_inst_569_dout;
wire [11:8] ram16sdp_inst_570_dout;
wire [15:12] ram16sdp_inst_571_dout;
wire [19:16] ram16sdp_inst_572_dout;
wire [23:20] ram16sdp_inst_573_dout;
wire [27:24] ram16sdp_inst_574_dout;
wire [31:28] ram16sdp_inst_575_dout;
wire [3:0] ram16sdp_inst_576_dout;
wire [7:4] ram16sdp_inst_577_dout;
wire [11:8] ram16sdp_inst_578_dout;
wire [15:12] ram16sdp_inst_579_dout;
wire [19:16] ram16sdp_inst_580_dout;
wire [23:20] ram16sdp_inst_581_dout;
wire [27:24] ram16sdp_inst_582_dout;
wire [31:28] ram16sdp_inst_583_dout;
wire [3:0] ram16sdp_inst_584_dout;
wire [7:4] ram16sdp_inst_585_dout;
wire [11:8] ram16sdp_inst_586_dout;
wire [15:12] ram16sdp_inst_587_dout;
wire [19:16] ram16sdp_inst_588_dout;
wire [23:20] ram16sdp_inst_589_dout;
wire [27:24] ram16sdp_inst_590_dout;
wire [31:28] ram16sdp_inst_591_dout;
wire [3:0] ram16sdp_inst_592_dout;
wire [7:4] ram16sdp_inst_593_dout;
wire [11:8] ram16sdp_inst_594_dout;
wire [15:12] ram16sdp_inst_595_dout;
wire [19:16] ram16sdp_inst_596_dout;
wire [23:20] ram16sdp_inst_597_dout;
wire [27:24] ram16sdp_inst_598_dout;
wire [31:28] ram16sdp_inst_599_dout;
wire [3:0] ram16sdp_inst_600_dout;
wire [7:4] ram16sdp_inst_601_dout;
wire [11:8] ram16sdp_inst_602_dout;
wire [15:12] ram16sdp_inst_603_dout;
wire [19:16] ram16sdp_inst_604_dout;
wire [23:20] ram16sdp_inst_605_dout;
wire [27:24] ram16sdp_inst_606_dout;
wire [31:28] ram16sdp_inst_607_dout;
wire [3:0] ram16sdp_inst_608_dout;
wire [7:4] ram16sdp_inst_609_dout;
wire [11:8] ram16sdp_inst_610_dout;
wire [15:12] ram16sdp_inst_611_dout;
wire [19:16] ram16sdp_inst_612_dout;
wire [23:20] ram16sdp_inst_613_dout;
wire [27:24] ram16sdp_inst_614_dout;
wire [31:28] ram16sdp_inst_615_dout;
wire [3:0] ram16sdp_inst_616_dout;
wire [7:4] ram16sdp_inst_617_dout;
wire [11:8] ram16sdp_inst_618_dout;
wire [15:12] ram16sdp_inst_619_dout;
wire [19:16] ram16sdp_inst_620_dout;
wire [23:20] ram16sdp_inst_621_dout;
wire [27:24] ram16sdp_inst_622_dout;
wire [31:28] ram16sdp_inst_623_dout;
wire [3:0] ram16sdp_inst_624_dout;
wire [7:4] ram16sdp_inst_625_dout;
wire [11:8] ram16sdp_inst_626_dout;
wire [15:12] ram16sdp_inst_627_dout;
wire [19:16] ram16sdp_inst_628_dout;
wire [23:20] ram16sdp_inst_629_dout;
wire [27:24] ram16sdp_inst_630_dout;
wire [31:28] ram16sdp_inst_631_dout;
wire [3:0] ram16sdp_inst_632_dout;
wire [7:4] ram16sdp_inst_633_dout;
wire [11:8] ram16sdp_inst_634_dout;
wire [15:12] ram16sdp_inst_635_dout;
wire [19:16] ram16sdp_inst_636_dout;
wire [23:20] ram16sdp_inst_637_dout;
wire [27:24] ram16sdp_inst_638_dout;
wire [31:28] ram16sdp_inst_639_dout;
wire [3:0] ram16sdp_inst_640_dout;
wire [7:4] ram16sdp_inst_641_dout;
wire [11:8] ram16sdp_inst_642_dout;
wire [15:12] ram16sdp_inst_643_dout;
wire [19:16] ram16sdp_inst_644_dout;
wire [23:20] ram16sdp_inst_645_dout;
wire [27:24] ram16sdp_inst_646_dout;
wire [31:28] ram16sdp_inst_647_dout;
wire [3:0] ram16sdp_inst_648_dout;
wire [7:4] ram16sdp_inst_649_dout;
wire [11:8] ram16sdp_inst_650_dout;
wire [15:12] ram16sdp_inst_651_dout;
wire [19:16] ram16sdp_inst_652_dout;
wire [23:20] ram16sdp_inst_653_dout;
wire [27:24] ram16sdp_inst_654_dout;
wire [31:28] ram16sdp_inst_655_dout;
wire [3:0] ram16sdp_inst_656_dout;
wire [7:4] ram16sdp_inst_657_dout;
wire [11:8] ram16sdp_inst_658_dout;
wire [15:12] ram16sdp_inst_659_dout;
wire [19:16] ram16sdp_inst_660_dout;
wire [23:20] ram16sdp_inst_661_dout;
wire [27:24] ram16sdp_inst_662_dout;
wire [31:28] ram16sdp_inst_663_dout;
wire [3:0] ram16sdp_inst_664_dout;
wire [7:4] ram16sdp_inst_665_dout;
wire [11:8] ram16sdp_inst_666_dout;
wire [15:12] ram16sdp_inst_667_dout;
wire [19:16] ram16sdp_inst_668_dout;
wire [23:20] ram16sdp_inst_669_dout;
wire [27:24] ram16sdp_inst_670_dout;
wire [31:28] ram16sdp_inst_671_dout;
wire [3:0] ram16sdp_inst_672_dout;
wire [7:4] ram16sdp_inst_673_dout;
wire [11:8] ram16sdp_inst_674_dout;
wire [15:12] ram16sdp_inst_675_dout;
wire [19:16] ram16sdp_inst_676_dout;
wire [23:20] ram16sdp_inst_677_dout;
wire [27:24] ram16sdp_inst_678_dout;
wire [31:28] ram16sdp_inst_679_dout;
wire [3:0] ram16sdp_inst_680_dout;
wire [7:4] ram16sdp_inst_681_dout;
wire [11:8] ram16sdp_inst_682_dout;
wire [15:12] ram16sdp_inst_683_dout;
wire [19:16] ram16sdp_inst_684_dout;
wire [23:20] ram16sdp_inst_685_dout;
wire [27:24] ram16sdp_inst_686_dout;
wire [31:28] ram16sdp_inst_687_dout;
wire [3:0] ram16sdp_inst_688_dout;
wire [7:4] ram16sdp_inst_689_dout;
wire [11:8] ram16sdp_inst_690_dout;
wire [15:12] ram16sdp_inst_691_dout;
wire [19:16] ram16sdp_inst_692_dout;
wire [23:20] ram16sdp_inst_693_dout;
wire [27:24] ram16sdp_inst_694_dout;
wire [31:28] ram16sdp_inst_695_dout;
wire [3:0] ram16sdp_inst_696_dout;
wire [7:4] ram16sdp_inst_697_dout;
wire [11:8] ram16sdp_inst_698_dout;
wire [15:12] ram16sdp_inst_699_dout;
wire [19:16] ram16sdp_inst_700_dout;
wire [23:20] ram16sdp_inst_701_dout;
wire [27:24] ram16sdp_inst_702_dout;
wire [31:28] ram16sdp_inst_703_dout;
wire [3:0] ram16sdp_inst_704_dout;
wire [7:4] ram16sdp_inst_705_dout;
wire [11:8] ram16sdp_inst_706_dout;
wire [15:12] ram16sdp_inst_707_dout;
wire [19:16] ram16sdp_inst_708_dout;
wire [23:20] ram16sdp_inst_709_dout;
wire [27:24] ram16sdp_inst_710_dout;
wire [31:28] ram16sdp_inst_711_dout;
wire [3:0] ram16sdp_inst_712_dout;
wire [7:4] ram16sdp_inst_713_dout;
wire [11:8] ram16sdp_inst_714_dout;
wire [15:12] ram16sdp_inst_715_dout;
wire [19:16] ram16sdp_inst_716_dout;
wire [23:20] ram16sdp_inst_717_dout;
wire [27:24] ram16sdp_inst_718_dout;
wire [31:28] ram16sdp_inst_719_dout;
wire [3:0] ram16sdp_inst_720_dout;
wire [7:4] ram16sdp_inst_721_dout;
wire [11:8] ram16sdp_inst_722_dout;
wire [15:12] ram16sdp_inst_723_dout;
wire [19:16] ram16sdp_inst_724_dout;
wire [23:20] ram16sdp_inst_725_dout;
wire [27:24] ram16sdp_inst_726_dout;
wire [31:28] ram16sdp_inst_727_dout;
wire [3:0] ram16sdp_inst_728_dout;
wire [7:4] ram16sdp_inst_729_dout;
wire [11:8] ram16sdp_inst_730_dout;
wire [15:12] ram16sdp_inst_731_dout;
wire [19:16] ram16sdp_inst_732_dout;
wire [23:20] ram16sdp_inst_733_dout;
wire [27:24] ram16sdp_inst_734_dout;
wire [31:28] ram16sdp_inst_735_dout;
wire [3:0] ram16sdp_inst_736_dout;
wire [7:4] ram16sdp_inst_737_dout;
wire [11:8] ram16sdp_inst_738_dout;
wire [15:12] ram16sdp_inst_739_dout;
wire [19:16] ram16sdp_inst_740_dout;
wire [23:20] ram16sdp_inst_741_dout;
wire [27:24] ram16sdp_inst_742_dout;
wire [31:28] ram16sdp_inst_743_dout;
wire [3:0] ram16sdp_inst_744_dout;
wire [7:4] ram16sdp_inst_745_dout;
wire [11:8] ram16sdp_inst_746_dout;
wire [15:12] ram16sdp_inst_747_dout;
wire [19:16] ram16sdp_inst_748_dout;
wire [23:20] ram16sdp_inst_749_dout;
wire [27:24] ram16sdp_inst_750_dout;
wire [31:28] ram16sdp_inst_751_dout;
wire [3:0] ram16sdp_inst_752_dout;
wire [7:4] ram16sdp_inst_753_dout;
wire [11:8] ram16sdp_inst_754_dout;
wire [15:12] ram16sdp_inst_755_dout;
wire [19:16] ram16sdp_inst_756_dout;
wire [23:20] ram16sdp_inst_757_dout;
wire [27:24] ram16sdp_inst_758_dout;
wire [31:28] ram16sdp_inst_759_dout;
wire [3:0] ram16sdp_inst_760_dout;
wire [7:4] ram16sdp_inst_761_dout;
wire [11:8] ram16sdp_inst_762_dout;
wire [15:12] ram16sdp_inst_763_dout;
wire [19:16] ram16sdp_inst_764_dout;
wire [23:20] ram16sdp_inst_765_dout;
wire [27:24] ram16sdp_inst_766_dout;
wire [31:28] ram16sdp_inst_767_dout;
wire [3:0] ram16sdp_inst_768_dout;
wire [7:4] ram16sdp_inst_769_dout;
wire [11:8] ram16sdp_inst_770_dout;
wire [15:12] ram16sdp_inst_771_dout;
wire [19:16] ram16sdp_inst_772_dout;
wire [23:20] ram16sdp_inst_773_dout;
wire [27:24] ram16sdp_inst_774_dout;
wire [31:28] ram16sdp_inst_775_dout;
wire [3:0] ram16sdp_inst_776_dout;
wire [7:4] ram16sdp_inst_777_dout;
wire [11:8] ram16sdp_inst_778_dout;
wire [15:12] ram16sdp_inst_779_dout;
wire [19:16] ram16sdp_inst_780_dout;
wire [23:20] ram16sdp_inst_781_dout;
wire [27:24] ram16sdp_inst_782_dout;
wire [31:28] ram16sdp_inst_783_dout;
wire [3:0] ram16sdp_inst_784_dout;
wire [7:4] ram16sdp_inst_785_dout;
wire [11:8] ram16sdp_inst_786_dout;
wire [15:12] ram16sdp_inst_787_dout;
wire [19:16] ram16sdp_inst_788_dout;
wire [23:20] ram16sdp_inst_789_dout;
wire [27:24] ram16sdp_inst_790_dout;
wire [31:28] ram16sdp_inst_791_dout;
wire [3:0] ram16sdp_inst_792_dout;
wire [7:4] ram16sdp_inst_793_dout;
wire [11:8] ram16sdp_inst_794_dout;
wire [15:12] ram16sdp_inst_795_dout;
wire [19:16] ram16sdp_inst_796_dout;
wire [23:20] ram16sdp_inst_797_dout;
wire [27:24] ram16sdp_inst_798_dout;
wire [31:28] ram16sdp_inst_799_dout;
wire [3:0] ram16sdp_inst_800_dout;
wire [7:4] ram16sdp_inst_801_dout;
wire [11:8] ram16sdp_inst_802_dout;
wire [15:12] ram16sdp_inst_803_dout;
wire [19:16] ram16sdp_inst_804_dout;
wire [23:20] ram16sdp_inst_805_dout;
wire [27:24] ram16sdp_inst_806_dout;
wire [31:28] ram16sdp_inst_807_dout;
wire [3:0] ram16sdp_inst_808_dout;
wire [7:4] ram16sdp_inst_809_dout;
wire [11:8] ram16sdp_inst_810_dout;
wire [15:12] ram16sdp_inst_811_dout;
wire [19:16] ram16sdp_inst_812_dout;
wire [23:20] ram16sdp_inst_813_dout;
wire [27:24] ram16sdp_inst_814_dout;
wire [31:28] ram16sdp_inst_815_dout;
wire [3:0] ram16sdp_inst_816_dout;
wire [7:4] ram16sdp_inst_817_dout;
wire [11:8] ram16sdp_inst_818_dout;
wire [15:12] ram16sdp_inst_819_dout;
wire [19:16] ram16sdp_inst_820_dout;
wire [23:20] ram16sdp_inst_821_dout;
wire [27:24] ram16sdp_inst_822_dout;
wire [31:28] ram16sdp_inst_823_dout;
wire [3:0] ram16sdp_inst_824_dout;
wire [7:4] ram16sdp_inst_825_dout;
wire [11:8] ram16sdp_inst_826_dout;
wire [15:12] ram16sdp_inst_827_dout;
wire [19:16] ram16sdp_inst_828_dout;
wire [23:20] ram16sdp_inst_829_dout;
wire [27:24] ram16sdp_inst_830_dout;
wire [31:28] ram16sdp_inst_831_dout;
wire [3:0] ram16sdp_inst_832_dout;
wire [7:4] ram16sdp_inst_833_dout;
wire [11:8] ram16sdp_inst_834_dout;
wire [15:12] ram16sdp_inst_835_dout;
wire [19:16] ram16sdp_inst_836_dout;
wire [23:20] ram16sdp_inst_837_dout;
wire [27:24] ram16sdp_inst_838_dout;
wire [31:28] ram16sdp_inst_839_dout;
wire [3:0] ram16sdp_inst_840_dout;
wire [7:4] ram16sdp_inst_841_dout;
wire [11:8] ram16sdp_inst_842_dout;
wire [15:12] ram16sdp_inst_843_dout;
wire [19:16] ram16sdp_inst_844_dout;
wire [23:20] ram16sdp_inst_845_dout;
wire [27:24] ram16sdp_inst_846_dout;
wire [31:28] ram16sdp_inst_847_dout;
wire [3:0] ram16sdp_inst_848_dout;
wire [7:4] ram16sdp_inst_849_dout;
wire [11:8] ram16sdp_inst_850_dout;
wire [15:12] ram16sdp_inst_851_dout;
wire [19:16] ram16sdp_inst_852_dout;
wire [23:20] ram16sdp_inst_853_dout;
wire [27:24] ram16sdp_inst_854_dout;
wire [31:28] ram16sdp_inst_855_dout;
wire [3:0] ram16sdp_inst_856_dout;
wire [7:4] ram16sdp_inst_857_dout;
wire [11:8] ram16sdp_inst_858_dout;
wire [15:12] ram16sdp_inst_859_dout;
wire [19:16] ram16sdp_inst_860_dout;
wire [23:20] ram16sdp_inst_861_dout;
wire [27:24] ram16sdp_inst_862_dout;
wire [31:28] ram16sdp_inst_863_dout;
wire [3:0] ram16sdp_inst_864_dout;
wire [7:4] ram16sdp_inst_865_dout;
wire [11:8] ram16sdp_inst_866_dout;
wire [15:12] ram16sdp_inst_867_dout;
wire [19:16] ram16sdp_inst_868_dout;
wire [23:20] ram16sdp_inst_869_dout;
wire [27:24] ram16sdp_inst_870_dout;
wire [31:28] ram16sdp_inst_871_dout;
wire [3:0] ram16sdp_inst_872_dout;
wire [7:4] ram16sdp_inst_873_dout;
wire [11:8] ram16sdp_inst_874_dout;
wire [15:12] ram16sdp_inst_875_dout;
wire [19:16] ram16sdp_inst_876_dout;
wire [23:20] ram16sdp_inst_877_dout;
wire [27:24] ram16sdp_inst_878_dout;
wire [31:28] ram16sdp_inst_879_dout;
wire [3:0] ram16sdp_inst_880_dout;
wire [7:4] ram16sdp_inst_881_dout;
wire [11:8] ram16sdp_inst_882_dout;
wire [15:12] ram16sdp_inst_883_dout;
wire [19:16] ram16sdp_inst_884_dout;
wire [23:20] ram16sdp_inst_885_dout;
wire [27:24] ram16sdp_inst_886_dout;
wire [31:28] ram16sdp_inst_887_dout;
wire [3:0] ram16sdp_inst_888_dout;
wire [7:4] ram16sdp_inst_889_dout;
wire [11:8] ram16sdp_inst_890_dout;
wire [15:12] ram16sdp_inst_891_dout;
wire [19:16] ram16sdp_inst_892_dout;
wire [23:20] ram16sdp_inst_893_dout;
wire [27:24] ram16sdp_inst_894_dout;
wire [31:28] ram16sdp_inst_895_dout;
wire [3:0] ram16sdp_inst_896_dout;
wire [7:4] ram16sdp_inst_897_dout;
wire [11:8] ram16sdp_inst_898_dout;
wire [15:12] ram16sdp_inst_899_dout;
wire [19:16] ram16sdp_inst_900_dout;
wire [23:20] ram16sdp_inst_901_dout;
wire [27:24] ram16sdp_inst_902_dout;
wire [31:28] ram16sdp_inst_903_dout;
wire [3:0] ram16sdp_inst_904_dout;
wire [7:4] ram16sdp_inst_905_dout;
wire [11:8] ram16sdp_inst_906_dout;
wire [15:12] ram16sdp_inst_907_dout;
wire [19:16] ram16sdp_inst_908_dout;
wire [23:20] ram16sdp_inst_909_dout;
wire [27:24] ram16sdp_inst_910_dout;
wire [31:28] ram16sdp_inst_911_dout;
wire [3:0] ram16sdp_inst_912_dout;
wire [7:4] ram16sdp_inst_913_dout;
wire [11:8] ram16sdp_inst_914_dout;
wire [15:12] ram16sdp_inst_915_dout;
wire [19:16] ram16sdp_inst_916_dout;
wire [23:20] ram16sdp_inst_917_dout;
wire [27:24] ram16sdp_inst_918_dout;
wire [31:28] ram16sdp_inst_919_dout;
wire [3:0] ram16sdp_inst_920_dout;
wire [7:4] ram16sdp_inst_921_dout;
wire [11:8] ram16sdp_inst_922_dout;
wire [15:12] ram16sdp_inst_923_dout;
wire [19:16] ram16sdp_inst_924_dout;
wire [23:20] ram16sdp_inst_925_dout;
wire [27:24] ram16sdp_inst_926_dout;
wire [31:28] ram16sdp_inst_927_dout;
wire [3:0] ram16sdp_inst_928_dout;
wire [7:4] ram16sdp_inst_929_dout;
wire [11:8] ram16sdp_inst_930_dout;
wire [15:12] ram16sdp_inst_931_dout;
wire [19:16] ram16sdp_inst_932_dout;
wire [23:20] ram16sdp_inst_933_dout;
wire [27:24] ram16sdp_inst_934_dout;
wire [31:28] ram16sdp_inst_935_dout;
wire [3:0] ram16sdp_inst_936_dout;
wire [7:4] ram16sdp_inst_937_dout;
wire [11:8] ram16sdp_inst_938_dout;
wire [15:12] ram16sdp_inst_939_dout;
wire [19:16] ram16sdp_inst_940_dout;
wire [23:20] ram16sdp_inst_941_dout;
wire [27:24] ram16sdp_inst_942_dout;
wire [31:28] ram16sdp_inst_943_dout;
wire [3:0] ram16sdp_inst_944_dout;
wire [7:4] ram16sdp_inst_945_dout;
wire [11:8] ram16sdp_inst_946_dout;
wire [15:12] ram16sdp_inst_947_dout;
wire [19:16] ram16sdp_inst_948_dout;
wire [23:20] ram16sdp_inst_949_dout;
wire [27:24] ram16sdp_inst_950_dout;
wire [31:28] ram16sdp_inst_951_dout;
wire [3:0] ram16sdp_inst_952_dout;
wire [7:4] ram16sdp_inst_953_dout;
wire [11:8] ram16sdp_inst_954_dout;
wire [15:12] ram16sdp_inst_955_dout;
wire [19:16] ram16sdp_inst_956_dout;
wire [23:20] ram16sdp_inst_957_dout;
wire [27:24] ram16sdp_inst_958_dout;
wire [31:28] ram16sdp_inst_959_dout;
wire [3:0] ram16sdp_inst_960_dout;
wire [7:4] ram16sdp_inst_961_dout;
wire [11:8] ram16sdp_inst_962_dout;
wire [15:12] ram16sdp_inst_963_dout;
wire [19:16] ram16sdp_inst_964_dout;
wire [23:20] ram16sdp_inst_965_dout;
wire [27:24] ram16sdp_inst_966_dout;
wire [31:28] ram16sdp_inst_967_dout;
wire [3:0] ram16sdp_inst_968_dout;
wire [7:4] ram16sdp_inst_969_dout;
wire [11:8] ram16sdp_inst_970_dout;
wire [15:12] ram16sdp_inst_971_dout;
wire [19:16] ram16sdp_inst_972_dout;
wire [23:20] ram16sdp_inst_973_dout;
wire [27:24] ram16sdp_inst_974_dout;
wire [31:28] ram16sdp_inst_975_dout;
wire [3:0] ram16sdp_inst_976_dout;
wire [7:4] ram16sdp_inst_977_dout;
wire [11:8] ram16sdp_inst_978_dout;
wire [15:12] ram16sdp_inst_979_dout;
wire [19:16] ram16sdp_inst_980_dout;
wire [23:20] ram16sdp_inst_981_dout;
wire [27:24] ram16sdp_inst_982_dout;
wire [31:28] ram16sdp_inst_983_dout;
wire [3:0] ram16sdp_inst_984_dout;
wire [7:4] ram16sdp_inst_985_dout;
wire [11:8] ram16sdp_inst_986_dout;
wire [15:12] ram16sdp_inst_987_dout;
wire [19:16] ram16sdp_inst_988_dout;
wire [23:20] ram16sdp_inst_989_dout;
wire [27:24] ram16sdp_inst_990_dout;
wire [31:28] ram16sdp_inst_991_dout;
wire [3:0] ram16sdp_inst_992_dout;
wire [7:4] ram16sdp_inst_993_dout;
wire [11:8] ram16sdp_inst_994_dout;
wire [15:12] ram16sdp_inst_995_dout;
wire [19:16] ram16sdp_inst_996_dout;
wire [23:20] ram16sdp_inst_997_dout;
wire [27:24] ram16sdp_inst_998_dout;
wire [31:28] ram16sdp_inst_999_dout;
wire [3:0] ram16sdp_inst_1000_dout;
wire [7:4] ram16sdp_inst_1001_dout;
wire [11:8] ram16sdp_inst_1002_dout;
wire [15:12] ram16sdp_inst_1003_dout;
wire [19:16] ram16sdp_inst_1004_dout;
wire [23:20] ram16sdp_inst_1005_dout;
wire [27:24] ram16sdp_inst_1006_dout;
wire [31:28] ram16sdp_inst_1007_dout;
wire [3:0] ram16sdp_inst_1008_dout;
wire [7:4] ram16sdp_inst_1009_dout;
wire [11:8] ram16sdp_inst_1010_dout;
wire [15:12] ram16sdp_inst_1011_dout;
wire [19:16] ram16sdp_inst_1012_dout;
wire [23:20] ram16sdp_inst_1013_dout;
wire [27:24] ram16sdp_inst_1014_dout;
wire [31:28] ram16sdp_inst_1015_dout;
wire [3:0] ram16sdp_inst_1016_dout;
wire [7:4] ram16sdp_inst_1017_dout;
wire [11:8] ram16sdp_inst_1018_dout;
wire [15:12] ram16sdp_inst_1019_dout;
wire [19:16] ram16sdp_inst_1020_dout;
wire [23:20] ram16sdp_inst_1021_dout;
wire [27:24] ram16sdp_inst_1022_dout;
wire [31:28] ram16sdp_inst_1023_dout;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_125;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_252;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_314;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_419;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_464;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_487;
wire mux_o_488;
wire mux_o_489;
wire mux_o_490;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_494;
wire mux_o_495;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_501;
wire mux_o_502;
wire mux_o_503;
wire mux_o_504;
wire mux_o_505;
wire mux_o_506;
wire mux_o_508;
wire mux_o_509;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_515;
wire mux_o_516;
wire mux_o_517;
wire mux_o_518;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_524;
wire mux_o_525;
wire mux_o_526;
wire mux_o_527;
wire mux_o_528;
wire mux_o_529;
wire mux_o_530;
wire mux_o_531;
wire mux_o_532;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_539;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_557;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_566;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_571;
wire mux_o_572;
wire mux_o_573;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_588;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_599;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_613;
wire mux_o_614;
wire mux_o_615;
wire mux_o_616;
wire mux_o_617;
wire mux_o_618;
wire mux_o_619;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_627;
wire mux_o_628;
wire mux_o_629;
wire mux_o_630;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_641;
wire mux_o_642;
wire mux_o_643;
wire mux_o_644;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_650;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_655;
wire mux_o_656;
wire mux_o_657;
wire mux_o_658;
wire mux_o_659;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_681;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_692;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_711;
wire mux_o_712;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_725;
wire mux_o_726;
wire mux_o_727;
wire mux_o_728;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_734;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_739;
wire mux_o_740;
wire mux_o_741;
wire mux_o_742;
wire mux_o_743;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_749;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_753;
wire mux_o_754;
wire mux_o_755;
wire mux_o_756;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_762;
wire mux_o_763;
wire mux_o_764;
wire mux_o_765;
wire mux_o_766;
wire mux_o_767;
wire mux_o_768;
wire mux_o_769;
wire mux_o_770;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_774;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_779;
wire mux_o_780;
wire mux_o_781;
wire mux_o_782;
wire mux_o_783;
wire mux_o_784;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_794;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_798;
wire mux_o_799;
wire mux_o_800;
wire mux_o_801;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_805;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_809;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_813;
wire mux_o_814;
wire mux_o_815;
wire mux_o_816;
wire mux_o_817;
wire mux_o_818;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_824;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_830;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_836;
wire mux_o_837;
wire mux_o_838;
wire mux_o_839;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_846;
wire mux_o_847;
wire mux_o_848;
wire mux_o_849;
wire mux_o_850;
wire mux_o_851;
wire mux_o_852;
wire mux_o_853;
wire mux_o_854;
wire mux_o_855;
wire mux_o_856;
wire mux_o_857;
wire mux_o_858;
wire mux_o_859;
wire mux_o_860;
wire mux_o_861;
wire mux_o_862;
wire mux_o_863;
wire mux_o_864;
wire mux_o_865;
wire mux_o_866;
wire mux_o_867;
wire mux_o_868;
wire mux_o_869;
wire mux_o_870;
wire mux_o_871;
wire mux_o_872;
wire mux_o_873;
wire mux_o_874;
wire mux_o_875;
wire mux_o_876;
wire mux_o_877;
wire mux_o_878;
wire mux_o_879;
wire mux_o_880;
wire mux_o_881;
wire mux_o_882;
wire mux_o_883;
wire mux_o_884;
wire mux_o_885;
wire mux_o_886;
wire mux_o_887;
wire mux_o_889;
wire mux_o_890;
wire mux_o_891;
wire mux_o_892;
wire mux_o_893;
wire mux_o_894;
wire mux_o_895;
wire mux_o_896;
wire mux_o_897;
wire mux_o_898;
wire mux_o_899;
wire mux_o_900;
wire mux_o_901;
wire mux_o_902;
wire mux_o_903;
wire mux_o_904;
wire mux_o_905;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_914;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_929;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_934;
wire mux_o_935;
wire mux_o_936;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_944;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_951;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire mux_o_959;
wire mux_o_960;
wire mux_o_961;
wire mux_o_962;
wire mux_o_963;
wire mux_o_964;
wire mux_o_965;
wire mux_o_966;
wire mux_o_967;
wire mux_o_968;
wire mux_o_969;
wire mux_o_970;
wire mux_o_971;
wire mux_o_972;
wire mux_o_973;
wire mux_o_974;
wire mux_o_975;
wire mux_o_976;
wire mux_o_977;
wire mux_o_978;
wire mux_o_979;
wire mux_o_980;
wire mux_o_981;
wire mux_o_982;
wire mux_o_983;
wire mux_o_984;
wire mux_o_985;
wire mux_o_986;
wire mux_o_987;
wire mux_o_988;
wire mux_o_989;
wire mux_o_990;
wire mux_o_991;
wire mux_o_992;
wire mux_o_993;
wire mux_o_994;
wire mux_o_995;
wire mux_o_996;
wire mux_o_997;
wire mux_o_998;
wire mux_o_999;
wire mux_o_1000;
wire mux_o_1001;
wire mux_o_1002;
wire mux_o_1003;
wire mux_o_1004;
wire mux_o_1005;
wire mux_o_1006;
wire mux_o_1007;
wire mux_o_1008;
wire mux_o_1009;
wire mux_o_1010;
wire mux_o_1011;
wire mux_o_1012;
wire mux_o_1013;
wire mux_o_1014;
wire mux_o_1016;
wire mux_o_1017;
wire mux_o_1018;
wire mux_o_1019;
wire mux_o_1020;
wire mux_o_1021;
wire mux_o_1022;
wire mux_o_1023;
wire mux_o_1024;
wire mux_o_1025;
wire mux_o_1026;
wire mux_o_1027;
wire mux_o_1028;
wire mux_o_1029;
wire mux_o_1030;
wire mux_o_1031;
wire mux_o_1032;
wire mux_o_1033;
wire mux_o_1034;
wire mux_o_1035;
wire mux_o_1036;
wire mux_o_1037;
wire mux_o_1038;
wire mux_o_1039;
wire mux_o_1040;
wire mux_o_1041;
wire mux_o_1042;
wire mux_o_1043;
wire mux_o_1044;
wire mux_o_1045;
wire mux_o_1046;
wire mux_o_1047;
wire mux_o_1048;
wire mux_o_1049;
wire mux_o_1050;
wire mux_o_1051;
wire mux_o_1052;
wire mux_o_1053;
wire mux_o_1054;
wire mux_o_1055;
wire mux_o_1056;
wire mux_o_1057;
wire mux_o_1058;
wire mux_o_1059;
wire mux_o_1060;
wire mux_o_1061;
wire mux_o_1062;
wire mux_o_1063;
wire mux_o_1064;
wire mux_o_1065;
wire mux_o_1066;
wire mux_o_1067;
wire mux_o_1068;
wire mux_o_1069;
wire mux_o_1070;
wire mux_o_1071;
wire mux_o_1072;
wire mux_o_1073;
wire mux_o_1074;
wire mux_o_1075;
wire mux_o_1076;
wire mux_o_1077;
wire mux_o_1078;
wire mux_o_1079;
wire mux_o_1080;
wire mux_o_1081;
wire mux_o_1082;
wire mux_o_1083;
wire mux_o_1084;
wire mux_o_1085;
wire mux_o_1086;
wire mux_o_1087;
wire mux_o_1088;
wire mux_o_1089;
wire mux_o_1090;
wire mux_o_1091;
wire mux_o_1092;
wire mux_o_1093;
wire mux_o_1094;
wire mux_o_1095;
wire mux_o_1096;
wire mux_o_1097;
wire mux_o_1098;
wire mux_o_1099;
wire mux_o_1100;
wire mux_o_1101;
wire mux_o_1102;
wire mux_o_1103;
wire mux_o_1104;
wire mux_o_1105;
wire mux_o_1106;
wire mux_o_1107;
wire mux_o_1108;
wire mux_o_1109;
wire mux_o_1110;
wire mux_o_1111;
wire mux_o_1112;
wire mux_o_1113;
wire mux_o_1114;
wire mux_o_1115;
wire mux_o_1116;
wire mux_o_1117;
wire mux_o_1118;
wire mux_o_1119;
wire mux_o_1120;
wire mux_o_1121;
wire mux_o_1122;
wire mux_o_1123;
wire mux_o_1124;
wire mux_o_1125;
wire mux_o_1126;
wire mux_o_1127;
wire mux_o_1128;
wire mux_o_1129;
wire mux_o_1130;
wire mux_o_1131;
wire mux_o_1132;
wire mux_o_1133;
wire mux_o_1134;
wire mux_o_1135;
wire mux_o_1136;
wire mux_o_1137;
wire mux_o_1138;
wire mux_o_1139;
wire mux_o_1140;
wire mux_o_1141;
wire mux_o_1143;
wire mux_o_1144;
wire mux_o_1145;
wire mux_o_1146;
wire mux_o_1147;
wire mux_o_1148;
wire mux_o_1149;
wire mux_o_1150;
wire mux_o_1151;
wire mux_o_1152;
wire mux_o_1153;
wire mux_o_1154;
wire mux_o_1155;
wire mux_o_1156;
wire mux_o_1157;
wire mux_o_1158;
wire mux_o_1159;
wire mux_o_1160;
wire mux_o_1161;
wire mux_o_1162;
wire mux_o_1163;
wire mux_o_1164;
wire mux_o_1165;
wire mux_o_1166;
wire mux_o_1167;
wire mux_o_1168;
wire mux_o_1169;
wire mux_o_1170;
wire mux_o_1171;
wire mux_o_1172;
wire mux_o_1173;
wire mux_o_1174;
wire mux_o_1175;
wire mux_o_1176;
wire mux_o_1177;
wire mux_o_1178;
wire mux_o_1179;
wire mux_o_1180;
wire mux_o_1181;
wire mux_o_1182;
wire mux_o_1183;
wire mux_o_1184;
wire mux_o_1185;
wire mux_o_1186;
wire mux_o_1187;
wire mux_o_1188;
wire mux_o_1189;
wire mux_o_1190;
wire mux_o_1191;
wire mux_o_1192;
wire mux_o_1193;
wire mux_o_1194;
wire mux_o_1195;
wire mux_o_1196;
wire mux_o_1197;
wire mux_o_1198;
wire mux_o_1199;
wire mux_o_1200;
wire mux_o_1201;
wire mux_o_1202;
wire mux_o_1203;
wire mux_o_1204;
wire mux_o_1205;
wire mux_o_1206;
wire mux_o_1207;
wire mux_o_1208;
wire mux_o_1209;
wire mux_o_1210;
wire mux_o_1211;
wire mux_o_1212;
wire mux_o_1213;
wire mux_o_1214;
wire mux_o_1215;
wire mux_o_1216;
wire mux_o_1217;
wire mux_o_1218;
wire mux_o_1219;
wire mux_o_1220;
wire mux_o_1221;
wire mux_o_1222;
wire mux_o_1223;
wire mux_o_1224;
wire mux_o_1225;
wire mux_o_1226;
wire mux_o_1227;
wire mux_o_1228;
wire mux_o_1229;
wire mux_o_1230;
wire mux_o_1231;
wire mux_o_1232;
wire mux_o_1233;
wire mux_o_1234;
wire mux_o_1235;
wire mux_o_1236;
wire mux_o_1237;
wire mux_o_1238;
wire mux_o_1239;
wire mux_o_1240;
wire mux_o_1241;
wire mux_o_1242;
wire mux_o_1243;
wire mux_o_1244;
wire mux_o_1245;
wire mux_o_1246;
wire mux_o_1247;
wire mux_o_1248;
wire mux_o_1249;
wire mux_o_1250;
wire mux_o_1251;
wire mux_o_1252;
wire mux_o_1253;
wire mux_o_1254;
wire mux_o_1255;
wire mux_o_1256;
wire mux_o_1257;
wire mux_o_1258;
wire mux_o_1259;
wire mux_o_1260;
wire mux_o_1261;
wire mux_o_1262;
wire mux_o_1263;
wire mux_o_1264;
wire mux_o_1265;
wire mux_o_1266;
wire mux_o_1267;
wire mux_o_1268;
wire mux_o_1270;
wire mux_o_1271;
wire mux_o_1272;
wire mux_o_1273;
wire mux_o_1274;
wire mux_o_1275;
wire mux_o_1276;
wire mux_o_1277;
wire mux_o_1278;
wire mux_o_1279;
wire mux_o_1280;
wire mux_o_1281;
wire mux_o_1282;
wire mux_o_1283;
wire mux_o_1284;
wire mux_o_1285;
wire mux_o_1286;
wire mux_o_1287;
wire mux_o_1288;
wire mux_o_1289;
wire mux_o_1290;
wire mux_o_1291;
wire mux_o_1292;
wire mux_o_1293;
wire mux_o_1294;
wire mux_o_1295;
wire mux_o_1296;
wire mux_o_1297;
wire mux_o_1298;
wire mux_o_1299;
wire mux_o_1300;
wire mux_o_1301;
wire mux_o_1302;
wire mux_o_1303;
wire mux_o_1304;
wire mux_o_1305;
wire mux_o_1306;
wire mux_o_1307;
wire mux_o_1308;
wire mux_o_1309;
wire mux_o_1310;
wire mux_o_1311;
wire mux_o_1312;
wire mux_o_1313;
wire mux_o_1314;
wire mux_o_1315;
wire mux_o_1316;
wire mux_o_1317;
wire mux_o_1318;
wire mux_o_1319;
wire mux_o_1320;
wire mux_o_1321;
wire mux_o_1322;
wire mux_o_1323;
wire mux_o_1324;
wire mux_o_1325;
wire mux_o_1326;
wire mux_o_1327;
wire mux_o_1328;
wire mux_o_1329;
wire mux_o_1330;
wire mux_o_1331;
wire mux_o_1332;
wire mux_o_1333;
wire mux_o_1334;
wire mux_o_1335;
wire mux_o_1336;
wire mux_o_1337;
wire mux_o_1338;
wire mux_o_1339;
wire mux_o_1340;
wire mux_o_1341;
wire mux_o_1342;
wire mux_o_1343;
wire mux_o_1344;
wire mux_o_1345;
wire mux_o_1346;
wire mux_o_1347;
wire mux_o_1348;
wire mux_o_1349;
wire mux_o_1350;
wire mux_o_1351;
wire mux_o_1352;
wire mux_o_1353;
wire mux_o_1354;
wire mux_o_1355;
wire mux_o_1356;
wire mux_o_1357;
wire mux_o_1358;
wire mux_o_1359;
wire mux_o_1360;
wire mux_o_1361;
wire mux_o_1362;
wire mux_o_1363;
wire mux_o_1364;
wire mux_o_1365;
wire mux_o_1366;
wire mux_o_1367;
wire mux_o_1368;
wire mux_o_1369;
wire mux_o_1370;
wire mux_o_1371;
wire mux_o_1372;
wire mux_o_1373;
wire mux_o_1374;
wire mux_o_1375;
wire mux_o_1376;
wire mux_o_1377;
wire mux_o_1378;
wire mux_o_1379;
wire mux_o_1380;
wire mux_o_1381;
wire mux_o_1382;
wire mux_o_1383;
wire mux_o_1384;
wire mux_o_1385;
wire mux_o_1386;
wire mux_o_1387;
wire mux_o_1388;
wire mux_o_1389;
wire mux_o_1390;
wire mux_o_1391;
wire mux_o_1392;
wire mux_o_1393;
wire mux_o_1394;
wire mux_o_1395;
wire mux_o_1397;
wire mux_o_1398;
wire mux_o_1399;
wire mux_o_1400;
wire mux_o_1401;
wire mux_o_1402;
wire mux_o_1403;
wire mux_o_1404;
wire mux_o_1405;
wire mux_o_1406;
wire mux_o_1407;
wire mux_o_1408;
wire mux_o_1409;
wire mux_o_1410;
wire mux_o_1411;
wire mux_o_1412;
wire mux_o_1413;
wire mux_o_1414;
wire mux_o_1415;
wire mux_o_1416;
wire mux_o_1417;
wire mux_o_1418;
wire mux_o_1419;
wire mux_o_1420;
wire mux_o_1421;
wire mux_o_1422;
wire mux_o_1423;
wire mux_o_1424;
wire mux_o_1425;
wire mux_o_1426;
wire mux_o_1427;
wire mux_o_1428;
wire mux_o_1429;
wire mux_o_1430;
wire mux_o_1431;
wire mux_o_1432;
wire mux_o_1433;
wire mux_o_1434;
wire mux_o_1435;
wire mux_o_1436;
wire mux_o_1437;
wire mux_o_1438;
wire mux_o_1439;
wire mux_o_1440;
wire mux_o_1441;
wire mux_o_1442;
wire mux_o_1443;
wire mux_o_1444;
wire mux_o_1445;
wire mux_o_1446;
wire mux_o_1447;
wire mux_o_1448;
wire mux_o_1449;
wire mux_o_1450;
wire mux_o_1451;
wire mux_o_1452;
wire mux_o_1453;
wire mux_o_1454;
wire mux_o_1455;
wire mux_o_1456;
wire mux_o_1457;
wire mux_o_1458;
wire mux_o_1459;
wire mux_o_1460;
wire mux_o_1461;
wire mux_o_1462;
wire mux_o_1463;
wire mux_o_1464;
wire mux_o_1465;
wire mux_o_1466;
wire mux_o_1467;
wire mux_o_1468;
wire mux_o_1469;
wire mux_o_1470;
wire mux_o_1471;
wire mux_o_1472;
wire mux_o_1473;
wire mux_o_1474;
wire mux_o_1475;
wire mux_o_1476;
wire mux_o_1477;
wire mux_o_1478;
wire mux_o_1479;
wire mux_o_1480;
wire mux_o_1481;
wire mux_o_1482;
wire mux_o_1483;
wire mux_o_1484;
wire mux_o_1485;
wire mux_o_1486;
wire mux_o_1487;
wire mux_o_1488;
wire mux_o_1489;
wire mux_o_1490;
wire mux_o_1491;
wire mux_o_1492;
wire mux_o_1493;
wire mux_o_1494;
wire mux_o_1495;
wire mux_o_1496;
wire mux_o_1497;
wire mux_o_1498;
wire mux_o_1499;
wire mux_o_1500;
wire mux_o_1501;
wire mux_o_1502;
wire mux_o_1503;
wire mux_o_1504;
wire mux_o_1505;
wire mux_o_1506;
wire mux_o_1507;
wire mux_o_1508;
wire mux_o_1509;
wire mux_o_1510;
wire mux_o_1511;
wire mux_o_1512;
wire mux_o_1513;
wire mux_o_1514;
wire mux_o_1515;
wire mux_o_1516;
wire mux_o_1517;
wire mux_o_1518;
wire mux_o_1519;
wire mux_o_1520;
wire mux_o_1521;
wire mux_o_1522;
wire mux_o_1524;
wire mux_o_1525;
wire mux_o_1526;
wire mux_o_1527;
wire mux_o_1528;
wire mux_o_1529;
wire mux_o_1530;
wire mux_o_1531;
wire mux_o_1532;
wire mux_o_1533;
wire mux_o_1534;
wire mux_o_1535;
wire mux_o_1536;
wire mux_o_1537;
wire mux_o_1538;
wire mux_o_1539;
wire mux_o_1540;
wire mux_o_1541;
wire mux_o_1542;
wire mux_o_1543;
wire mux_o_1544;
wire mux_o_1545;
wire mux_o_1546;
wire mux_o_1547;
wire mux_o_1548;
wire mux_o_1549;
wire mux_o_1550;
wire mux_o_1551;
wire mux_o_1552;
wire mux_o_1553;
wire mux_o_1554;
wire mux_o_1555;
wire mux_o_1556;
wire mux_o_1557;
wire mux_o_1558;
wire mux_o_1559;
wire mux_o_1560;
wire mux_o_1561;
wire mux_o_1562;
wire mux_o_1563;
wire mux_o_1564;
wire mux_o_1565;
wire mux_o_1566;
wire mux_o_1567;
wire mux_o_1568;
wire mux_o_1569;
wire mux_o_1570;
wire mux_o_1571;
wire mux_o_1572;
wire mux_o_1573;
wire mux_o_1574;
wire mux_o_1575;
wire mux_o_1576;
wire mux_o_1577;
wire mux_o_1578;
wire mux_o_1579;
wire mux_o_1580;
wire mux_o_1581;
wire mux_o_1582;
wire mux_o_1583;
wire mux_o_1584;
wire mux_o_1585;
wire mux_o_1586;
wire mux_o_1587;
wire mux_o_1588;
wire mux_o_1589;
wire mux_o_1590;
wire mux_o_1591;
wire mux_o_1592;
wire mux_o_1593;
wire mux_o_1594;
wire mux_o_1595;
wire mux_o_1596;
wire mux_o_1597;
wire mux_o_1598;
wire mux_o_1599;
wire mux_o_1600;
wire mux_o_1601;
wire mux_o_1602;
wire mux_o_1603;
wire mux_o_1604;
wire mux_o_1605;
wire mux_o_1606;
wire mux_o_1607;
wire mux_o_1608;
wire mux_o_1609;
wire mux_o_1610;
wire mux_o_1611;
wire mux_o_1612;
wire mux_o_1613;
wire mux_o_1614;
wire mux_o_1615;
wire mux_o_1616;
wire mux_o_1617;
wire mux_o_1618;
wire mux_o_1619;
wire mux_o_1620;
wire mux_o_1621;
wire mux_o_1622;
wire mux_o_1623;
wire mux_o_1624;
wire mux_o_1625;
wire mux_o_1626;
wire mux_o_1627;
wire mux_o_1628;
wire mux_o_1629;
wire mux_o_1630;
wire mux_o_1631;
wire mux_o_1632;
wire mux_o_1633;
wire mux_o_1634;
wire mux_o_1635;
wire mux_o_1636;
wire mux_o_1637;
wire mux_o_1638;
wire mux_o_1639;
wire mux_o_1640;
wire mux_o_1641;
wire mux_o_1642;
wire mux_o_1643;
wire mux_o_1644;
wire mux_o_1645;
wire mux_o_1646;
wire mux_o_1647;
wire mux_o_1648;
wire mux_o_1649;
wire mux_o_1651;
wire mux_o_1652;
wire mux_o_1653;
wire mux_o_1654;
wire mux_o_1655;
wire mux_o_1656;
wire mux_o_1657;
wire mux_o_1658;
wire mux_o_1659;
wire mux_o_1660;
wire mux_o_1661;
wire mux_o_1662;
wire mux_o_1663;
wire mux_o_1664;
wire mux_o_1665;
wire mux_o_1666;
wire mux_o_1667;
wire mux_o_1668;
wire mux_o_1669;
wire mux_o_1670;
wire mux_o_1671;
wire mux_o_1672;
wire mux_o_1673;
wire mux_o_1674;
wire mux_o_1675;
wire mux_o_1676;
wire mux_o_1677;
wire mux_o_1678;
wire mux_o_1679;
wire mux_o_1680;
wire mux_o_1681;
wire mux_o_1682;
wire mux_o_1683;
wire mux_o_1684;
wire mux_o_1685;
wire mux_o_1686;
wire mux_o_1687;
wire mux_o_1688;
wire mux_o_1689;
wire mux_o_1690;
wire mux_o_1691;
wire mux_o_1692;
wire mux_o_1693;
wire mux_o_1694;
wire mux_o_1695;
wire mux_o_1696;
wire mux_o_1697;
wire mux_o_1698;
wire mux_o_1699;
wire mux_o_1700;
wire mux_o_1701;
wire mux_o_1702;
wire mux_o_1703;
wire mux_o_1704;
wire mux_o_1705;
wire mux_o_1706;
wire mux_o_1707;
wire mux_o_1708;
wire mux_o_1709;
wire mux_o_1710;
wire mux_o_1711;
wire mux_o_1712;
wire mux_o_1713;
wire mux_o_1714;
wire mux_o_1715;
wire mux_o_1716;
wire mux_o_1717;
wire mux_o_1718;
wire mux_o_1719;
wire mux_o_1720;
wire mux_o_1721;
wire mux_o_1722;
wire mux_o_1723;
wire mux_o_1724;
wire mux_o_1725;
wire mux_o_1726;
wire mux_o_1727;
wire mux_o_1728;
wire mux_o_1729;
wire mux_o_1730;
wire mux_o_1731;
wire mux_o_1732;
wire mux_o_1733;
wire mux_o_1734;
wire mux_o_1735;
wire mux_o_1736;
wire mux_o_1737;
wire mux_o_1738;
wire mux_o_1739;
wire mux_o_1740;
wire mux_o_1741;
wire mux_o_1742;
wire mux_o_1743;
wire mux_o_1744;
wire mux_o_1745;
wire mux_o_1746;
wire mux_o_1747;
wire mux_o_1748;
wire mux_o_1749;
wire mux_o_1750;
wire mux_o_1751;
wire mux_o_1752;
wire mux_o_1753;
wire mux_o_1754;
wire mux_o_1755;
wire mux_o_1756;
wire mux_o_1757;
wire mux_o_1758;
wire mux_o_1759;
wire mux_o_1760;
wire mux_o_1761;
wire mux_o_1762;
wire mux_o_1763;
wire mux_o_1764;
wire mux_o_1765;
wire mux_o_1766;
wire mux_o_1767;
wire mux_o_1768;
wire mux_o_1769;
wire mux_o_1770;
wire mux_o_1771;
wire mux_o_1772;
wire mux_o_1773;
wire mux_o_1774;
wire mux_o_1775;
wire mux_o_1776;
wire mux_o_1778;
wire mux_o_1779;
wire mux_o_1780;
wire mux_o_1781;
wire mux_o_1782;
wire mux_o_1783;
wire mux_o_1784;
wire mux_o_1785;
wire mux_o_1786;
wire mux_o_1787;
wire mux_o_1788;
wire mux_o_1789;
wire mux_o_1790;
wire mux_o_1791;
wire mux_o_1792;
wire mux_o_1793;
wire mux_o_1794;
wire mux_o_1795;
wire mux_o_1796;
wire mux_o_1797;
wire mux_o_1798;
wire mux_o_1799;
wire mux_o_1800;
wire mux_o_1801;
wire mux_o_1802;
wire mux_o_1803;
wire mux_o_1804;
wire mux_o_1805;
wire mux_o_1806;
wire mux_o_1807;
wire mux_o_1808;
wire mux_o_1809;
wire mux_o_1810;
wire mux_o_1811;
wire mux_o_1812;
wire mux_o_1813;
wire mux_o_1814;
wire mux_o_1815;
wire mux_o_1816;
wire mux_o_1817;
wire mux_o_1818;
wire mux_o_1819;
wire mux_o_1820;
wire mux_o_1821;
wire mux_o_1822;
wire mux_o_1823;
wire mux_o_1824;
wire mux_o_1825;
wire mux_o_1826;
wire mux_o_1827;
wire mux_o_1828;
wire mux_o_1829;
wire mux_o_1830;
wire mux_o_1831;
wire mux_o_1832;
wire mux_o_1833;
wire mux_o_1834;
wire mux_o_1835;
wire mux_o_1836;
wire mux_o_1837;
wire mux_o_1838;
wire mux_o_1839;
wire mux_o_1840;
wire mux_o_1841;
wire mux_o_1842;
wire mux_o_1843;
wire mux_o_1844;
wire mux_o_1845;
wire mux_o_1846;
wire mux_o_1847;
wire mux_o_1848;
wire mux_o_1849;
wire mux_o_1850;
wire mux_o_1851;
wire mux_o_1852;
wire mux_o_1853;
wire mux_o_1854;
wire mux_o_1855;
wire mux_o_1856;
wire mux_o_1857;
wire mux_o_1858;
wire mux_o_1859;
wire mux_o_1860;
wire mux_o_1861;
wire mux_o_1862;
wire mux_o_1863;
wire mux_o_1864;
wire mux_o_1865;
wire mux_o_1866;
wire mux_o_1867;
wire mux_o_1868;
wire mux_o_1869;
wire mux_o_1870;
wire mux_o_1871;
wire mux_o_1872;
wire mux_o_1873;
wire mux_o_1874;
wire mux_o_1875;
wire mux_o_1876;
wire mux_o_1877;
wire mux_o_1878;
wire mux_o_1879;
wire mux_o_1880;
wire mux_o_1881;
wire mux_o_1882;
wire mux_o_1883;
wire mux_o_1884;
wire mux_o_1885;
wire mux_o_1886;
wire mux_o_1887;
wire mux_o_1888;
wire mux_o_1889;
wire mux_o_1890;
wire mux_o_1891;
wire mux_o_1892;
wire mux_o_1893;
wire mux_o_1894;
wire mux_o_1895;
wire mux_o_1896;
wire mux_o_1897;
wire mux_o_1898;
wire mux_o_1899;
wire mux_o_1900;
wire mux_o_1901;
wire mux_o_1902;
wire mux_o_1903;
wire mux_o_1905;
wire mux_o_1906;
wire mux_o_1907;
wire mux_o_1908;
wire mux_o_1909;
wire mux_o_1910;
wire mux_o_1911;
wire mux_o_1912;
wire mux_o_1913;
wire mux_o_1914;
wire mux_o_1915;
wire mux_o_1916;
wire mux_o_1917;
wire mux_o_1918;
wire mux_o_1919;
wire mux_o_1920;
wire mux_o_1921;
wire mux_o_1922;
wire mux_o_1923;
wire mux_o_1924;
wire mux_o_1925;
wire mux_o_1926;
wire mux_o_1927;
wire mux_o_1928;
wire mux_o_1929;
wire mux_o_1930;
wire mux_o_1931;
wire mux_o_1932;
wire mux_o_1933;
wire mux_o_1934;
wire mux_o_1935;
wire mux_o_1936;
wire mux_o_1937;
wire mux_o_1938;
wire mux_o_1939;
wire mux_o_1940;
wire mux_o_1941;
wire mux_o_1942;
wire mux_o_1943;
wire mux_o_1944;
wire mux_o_1945;
wire mux_o_1946;
wire mux_o_1947;
wire mux_o_1948;
wire mux_o_1949;
wire mux_o_1950;
wire mux_o_1951;
wire mux_o_1952;
wire mux_o_1953;
wire mux_o_1954;
wire mux_o_1955;
wire mux_o_1956;
wire mux_o_1957;
wire mux_o_1958;
wire mux_o_1959;
wire mux_o_1960;
wire mux_o_1961;
wire mux_o_1962;
wire mux_o_1963;
wire mux_o_1964;
wire mux_o_1965;
wire mux_o_1966;
wire mux_o_1967;
wire mux_o_1968;
wire mux_o_1969;
wire mux_o_1970;
wire mux_o_1971;
wire mux_o_1972;
wire mux_o_1973;
wire mux_o_1974;
wire mux_o_1975;
wire mux_o_1976;
wire mux_o_1977;
wire mux_o_1978;
wire mux_o_1979;
wire mux_o_1980;
wire mux_o_1981;
wire mux_o_1982;
wire mux_o_1983;
wire mux_o_1984;
wire mux_o_1985;
wire mux_o_1986;
wire mux_o_1987;
wire mux_o_1988;
wire mux_o_1989;
wire mux_o_1990;
wire mux_o_1991;
wire mux_o_1992;
wire mux_o_1993;
wire mux_o_1994;
wire mux_o_1995;
wire mux_o_1996;
wire mux_o_1997;
wire mux_o_1998;
wire mux_o_1999;
wire mux_o_2000;
wire mux_o_2001;
wire mux_o_2002;
wire mux_o_2003;
wire mux_o_2004;
wire mux_o_2005;
wire mux_o_2006;
wire mux_o_2007;
wire mux_o_2008;
wire mux_o_2009;
wire mux_o_2010;
wire mux_o_2011;
wire mux_o_2012;
wire mux_o_2013;
wire mux_o_2014;
wire mux_o_2015;
wire mux_o_2016;
wire mux_o_2017;
wire mux_o_2018;
wire mux_o_2019;
wire mux_o_2020;
wire mux_o_2021;
wire mux_o_2022;
wire mux_o_2023;
wire mux_o_2024;
wire mux_o_2025;
wire mux_o_2026;
wire mux_o_2027;
wire mux_o_2028;
wire mux_o_2029;
wire mux_o_2030;
wire mux_o_2032;
wire mux_o_2033;
wire mux_o_2034;
wire mux_o_2035;
wire mux_o_2036;
wire mux_o_2037;
wire mux_o_2038;
wire mux_o_2039;
wire mux_o_2040;
wire mux_o_2041;
wire mux_o_2042;
wire mux_o_2043;
wire mux_o_2044;
wire mux_o_2045;
wire mux_o_2046;
wire mux_o_2047;
wire mux_o_2048;
wire mux_o_2049;
wire mux_o_2050;
wire mux_o_2051;
wire mux_o_2052;
wire mux_o_2053;
wire mux_o_2054;
wire mux_o_2055;
wire mux_o_2056;
wire mux_o_2057;
wire mux_o_2058;
wire mux_o_2059;
wire mux_o_2060;
wire mux_o_2061;
wire mux_o_2062;
wire mux_o_2063;
wire mux_o_2064;
wire mux_o_2065;
wire mux_o_2066;
wire mux_o_2067;
wire mux_o_2068;
wire mux_o_2069;
wire mux_o_2070;
wire mux_o_2071;
wire mux_o_2072;
wire mux_o_2073;
wire mux_o_2074;
wire mux_o_2075;
wire mux_o_2076;
wire mux_o_2077;
wire mux_o_2078;
wire mux_o_2079;
wire mux_o_2080;
wire mux_o_2081;
wire mux_o_2082;
wire mux_o_2083;
wire mux_o_2084;
wire mux_o_2085;
wire mux_o_2086;
wire mux_o_2087;
wire mux_o_2088;
wire mux_o_2089;
wire mux_o_2090;
wire mux_o_2091;
wire mux_o_2092;
wire mux_o_2093;
wire mux_o_2094;
wire mux_o_2095;
wire mux_o_2096;
wire mux_o_2097;
wire mux_o_2098;
wire mux_o_2099;
wire mux_o_2100;
wire mux_o_2101;
wire mux_o_2102;
wire mux_o_2103;
wire mux_o_2104;
wire mux_o_2105;
wire mux_o_2106;
wire mux_o_2107;
wire mux_o_2108;
wire mux_o_2109;
wire mux_o_2110;
wire mux_o_2111;
wire mux_o_2112;
wire mux_o_2113;
wire mux_o_2114;
wire mux_o_2115;
wire mux_o_2116;
wire mux_o_2117;
wire mux_o_2118;
wire mux_o_2119;
wire mux_o_2120;
wire mux_o_2121;
wire mux_o_2122;
wire mux_o_2123;
wire mux_o_2124;
wire mux_o_2125;
wire mux_o_2126;
wire mux_o_2127;
wire mux_o_2128;
wire mux_o_2129;
wire mux_o_2130;
wire mux_o_2131;
wire mux_o_2132;
wire mux_o_2133;
wire mux_o_2134;
wire mux_o_2135;
wire mux_o_2136;
wire mux_o_2137;
wire mux_o_2138;
wire mux_o_2139;
wire mux_o_2140;
wire mux_o_2141;
wire mux_o_2142;
wire mux_o_2143;
wire mux_o_2144;
wire mux_o_2145;
wire mux_o_2146;
wire mux_o_2147;
wire mux_o_2148;
wire mux_o_2149;
wire mux_o_2150;
wire mux_o_2151;
wire mux_o_2152;
wire mux_o_2153;
wire mux_o_2154;
wire mux_o_2155;
wire mux_o_2156;
wire mux_o_2157;
wire mux_o_2159;
wire mux_o_2160;
wire mux_o_2161;
wire mux_o_2162;
wire mux_o_2163;
wire mux_o_2164;
wire mux_o_2165;
wire mux_o_2166;
wire mux_o_2167;
wire mux_o_2168;
wire mux_o_2169;
wire mux_o_2170;
wire mux_o_2171;
wire mux_o_2172;
wire mux_o_2173;
wire mux_o_2174;
wire mux_o_2175;
wire mux_o_2176;
wire mux_o_2177;
wire mux_o_2178;
wire mux_o_2179;
wire mux_o_2180;
wire mux_o_2181;
wire mux_o_2182;
wire mux_o_2183;
wire mux_o_2184;
wire mux_o_2185;
wire mux_o_2186;
wire mux_o_2187;
wire mux_o_2188;
wire mux_o_2189;
wire mux_o_2190;
wire mux_o_2191;
wire mux_o_2192;
wire mux_o_2193;
wire mux_o_2194;
wire mux_o_2195;
wire mux_o_2196;
wire mux_o_2197;
wire mux_o_2198;
wire mux_o_2199;
wire mux_o_2200;
wire mux_o_2201;
wire mux_o_2202;
wire mux_o_2203;
wire mux_o_2204;
wire mux_o_2205;
wire mux_o_2206;
wire mux_o_2207;
wire mux_o_2208;
wire mux_o_2209;
wire mux_o_2210;
wire mux_o_2211;
wire mux_o_2212;
wire mux_o_2213;
wire mux_o_2214;
wire mux_o_2215;
wire mux_o_2216;
wire mux_o_2217;
wire mux_o_2218;
wire mux_o_2219;
wire mux_o_2220;
wire mux_o_2221;
wire mux_o_2222;
wire mux_o_2223;
wire mux_o_2224;
wire mux_o_2225;
wire mux_o_2226;
wire mux_o_2227;
wire mux_o_2228;
wire mux_o_2229;
wire mux_o_2230;
wire mux_o_2231;
wire mux_o_2232;
wire mux_o_2233;
wire mux_o_2234;
wire mux_o_2235;
wire mux_o_2236;
wire mux_o_2237;
wire mux_o_2238;
wire mux_o_2239;
wire mux_o_2240;
wire mux_o_2241;
wire mux_o_2242;
wire mux_o_2243;
wire mux_o_2244;
wire mux_o_2245;
wire mux_o_2246;
wire mux_o_2247;
wire mux_o_2248;
wire mux_o_2249;
wire mux_o_2250;
wire mux_o_2251;
wire mux_o_2252;
wire mux_o_2253;
wire mux_o_2254;
wire mux_o_2255;
wire mux_o_2256;
wire mux_o_2257;
wire mux_o_2258;
wire mux_o_2259;
wire mux_o_2260;
wire mux_o_2261;
wire mux_o_2262;
wire mux_o_2263;
wire mux_o_2264;
wire mux_o_2265;
wire mux_o_2266;
wire mux_o_2267;
wire mux_o_2268;
wire mux_o_2269;
wire mux_o_2270;
wire mux_o_2271;
wire mux_o_2272;
wire mux_o_2273;
wire mux_o_2274;
wire mux_o_2275;
wire mux_o_2276;
wire mux_o_2277;
wire mux_o_2278;
wire mux_o_2279;
wire mux_o_2280;
wire mux_o_2281;
wire mux_o_2282;
wire mux_o_2283;
wire mux_o_2284;
wire mux_o_2286;
wire mux_o_2287;
wire mux_o_2288;
wire mux_o_2289;
wire mux_o_2290;
wire mux_o_2291;
wire mux_o_2292;
wire mux_o_2293;
wire mux_o_2294;
wire mux_o_2295;
wire mux_o_2296;
wire mux_o_2297;
wire mux_o_2298;
wire mux_o_2299;
wire mux_o_2300;
wire mux_o_2301;
wire mux_o_2302;
wire mux_o_2303;
wire mux_o_2304;
wire mux_o_2305;
wire mux_o_2306;
wire mux_o_2307;
wire mux_o_2308;
wire mux_o_2309;
wire mux_o_2310;
wire mux_o_2311;
wire mux_o_2312;
wire mux_o_2313;
wire mux_o_2314;
wire mux_o_2315;
wire mux_o_2316;
wire mux_o_2317;
wire mux_o_2318;
wire mux_o_2319;
wire mux_o_2320;
wire mux_o_2321;
wire mux_o_2322;
wire mux_o_2323;
wire mux_o_2324;
wire mux_o_2325;
wire mux_o_2326;
wire mux_o_2327;
wire mux_o_2328;
wire mux_o_2329;
wire mux_o_2330;
wire mux_o_2331;
wire mux_o_2332;
wire mux_o_2333;
wire mux_o_2334;
wire mux_o_2335;
wire mux_o_2336;
wire mux_o_2337;
wire mux_o_2338;
wire mux_o_2339;
wire mux_o_2340;
wire mux_o_2341;
wire mux_o_2342;
wire mux_o_2343;
wire mux_o_2344;
wire mux_o_2345;
wire mux_o_2346;
wire mux_o_2347;
wire mux_o_2348;
wire mux_o_2349;
wire mux_o_2350;
wire mux_o_2351;
wire mux_o_2352;
wire mux_o_2353;
wire mux_o_2354;
wire mux_o_2355;
wire mux_o_2356;
wire mux_o_2357;
wire mux_o_2358;
wire mux_o_2359;
wire mux_o_2360;
wire mux_o_2361;
wire mux_o_2362;
wire mux_o_2363;
wire mux_o_2364;
wire mux_o_2365;
wire mux_o_2366;
wire mux_o_2367;
wire mux_o_2368;
wire mux_o_2369;
wire mux_o_2370;
wire mux_o_2371;
wire mux_o_2372;
wire mux_o_2373;
wire mux_o_2374;
wire mux_o_2375;
wire mux_o_2376;
wire mux_o_2377;
wire mux_o_2378;
wire mux_o_2379;
wire mux_o_2380;
wire mux_o_2381;
wire mux_o_2382;
wire mux_o_2383;
wire mux_o_2384;
wire mux_o_2385;
wire mux_o_2386;
wire mux_o_2387;
wire mux_o_2388;
wire mux_o_2389;
wire mux_o_2390;
wire mux_o_2391;
wire mux_o_2392;
wire mux_o_2393;
wire mux_o_2394;
wire mux_o_2395;
wire mux_o_2396;
wire mux_o_2397;
wire mux_o_2398;
wire mux_o_2399;
wire mux_o_2400;
wire mux_o_2401;
wire mux_o_2402;
wire mux_o_2403;
wire mux_o_2404;
wire mux_o_2405;
wire mux_o_2406;
wire mux_o_2407;
wire mux_o_2408;
wire mux_o_2409;
wire mux_o_2410;
wire mux_o_2411;
wire mux_o_2413;
wire mux_o_2414;
wire mux_o_2415;
wire mux_o_2416;
wire mux_o_2417;
wire mux_o_2418;
wire mux_o_2419;
wire mux_o_2420;
wire mux_o_2421;
wire mux_o_2422;
wire mux_o_2423;
wire mux_o_2424;
wire mux_o_2425;
wire mux_o_2426;
wire mux_o_2427;
wire mux_o_2428;
wire mux_o_2429;
wire mux_o_2430;
wire mux_o_2431;
wire mux_o_2432;
wire mux_o_2433;
wire mux_o_2434;
wire mux_o_2435;
wire mux_o_2436;
wire mux_o_2437;
wire mux_o_2438;
wire mux_o_2439;
wire mux_o_2440;
wire mux_o_2441;
wire mux_o_2442;
wire mux_o_2443;
wire mux_o_2444;
wire mux_o_2445;
wire mux_o_2446;
wire mux_o_2447;
wire mux_o_2448;
wire mux_o_2449;
wire mux_o_2450;
wire mux_o_2451;
wire mux_o_2452;
wire mux_o_2453;
wire mux_o_2454;
wire mux_o_2455;
wire mux_o_2456;
wire mux_o_2457;
wire mux_o_2458;
wire mux_o_2459;
wire mux_o_2460;
wire mux_o_2461;
wire mux_o_2462;
wire mux_o_2463;
wire mux_o_2464;
wire mux_o_2465;
wire mux_o_2466;
wire mux_o_2467;
wire mux_o_2468;
wire mux_o_2469;
wire mux_o_2470;
wire mux_o_2471;
wire mux_o_2472;
wire mux_o_2473;
wire mux_o_2474;
wire mux_o_2475;
wire mux_o_2476;
wire mux_o_2477;
wire mux_o_2478;
wire mux_o_2479;
wire mux_o_2480;
wire mux_o_2481;
wire mux_o_2482;
wire mux_o_2483;
wire mux_o_2484;
wire mux_o_2485;
wire mux_o_2486;
wire mux_o_2487;
wire mux_o_2488;
wire mux_o_2489;
wire mux_o_2490;
wire mux_o_2491;
wire mux_o_2492;
wire mux_o_2493;
wire mux_o_2494;
wire mux_o_2495;
wire mux_o_2496;
wire mux_o_2497;
wire mux_o_2498;
wire mux_o_2499;
wire mux_o_2500;
wire mux_o_2501;
wire mux_o_2502;
wire mux_o_2503;
wire mux_o_2504;
wire mux_o_2505;
wire mux_o_2506;
wire mux_o_2507;
wire mux_o_2508;
wire mux_o_2509;
wire mux_o_2510;
wire mux_o_2511;
wire mux_o_2512;
wire mux_o_2513;
wire mux_o_2514;
wire mux_o_2515;
wire mux_o_2516;
wire mux_o_2517;
wire mux_o_2518;
wire mux_o_2519;
wire mux_o_2520;
wire mux_o_2521;
wire mux_o_2522;
wire mux_o_2523;
wire mux_o_2524;
wire mux_o_2525;
wire mux_o_2526;
wire mux_o_2527;
wire mux_o_2528;
wire mux_o_2529;
wire mux_o_2530;
wire mux_o_2531;
wire mux_o_2532;
wire mux_o_2533;
wire mux_o_2534;
wire mux_o_2535;
wire mux_o_2536;
wire mux_o_2537;
wire mux_o_2538;
wire mux_o_2540;
wire mux_o_2541;
wire mux_o_2542;
wire mux_o_2543;
wire mux_o_2544;
wire mux_o_2545;
wire mux_o_2546;
wire mux_o_2547;
wire mux_o_2548;
wire mux_o_2549;
wire mux_o_2550;
wire mux_o_2551;
wire mux_o_2552;
wire mux_o_2553;
wire mux_o_2554;
wire mux_o_2555;
wire mux_o_2556;
wire mux_o_2557;
wire mux_o_2558;
wire mux_o_2559;
wire mux_o_2560;
wire mux_o_2561;
wire mux_o_2562;
wire mux_o_2563;
wire mux_o_2564;
wire mux_o_2565;
wire mux_o_2566;
wire mux_o_2567;
wire mux_o_2568;
wire mux_o_2569;
wire mux_o_2570;
wire mux_o_2571;
wire mux_o_2572;
wire mux_o_2573;
wire mux_o_2574;
wire mux_o_2575;
wire mux_o_2576;
wire mux_o_2577;
wire mux_o_2578;
wire mux_o_2579;
wire mux_o_2580;
wire mux_o_2581;
wire mux_o_2582;
wire mux_o_2583;
wire mux_o_2584;
wire mux_o_2585;
wire mux_o_2586;
wire mux_o_2587;
wire mux_o_2588;
wire mux_o_2589;
wire mux_o_2590;
wire mux_o_2591;
wire mux_o_2592;
wire mux_o_2593;
wire mux_o_2594;
wire mux_o_2595;
wire mux_o_2596;
wire mux_o_2597;
wire mux_o_2598;
wire mux_o_2599;
wire mux_o_2600;
wire mux_o_2601;
wire mux_o_2602;
wire mux_o_2603;
wire mux_o_2604;
wire mux_o_2605;
wire mux_o_2606;
wire mux_o_2607;
wire mux_o_2608;
wire mux_o_2609;
wire mux_o_2610;
wire mux_o_2611;
wire mux_o_2612;
wire mux_o_2613;
wire mux_o_2614;
wire mux_o_2615;
wire mux_o_2616;
wire mux_o_2617;
wire mux_o_2618;
wire mux_o_2619;
wire mux_o_2620;
wire mux_o_2621;
wire mux_o_2622;
wire mux_o_2623;
wire mux_o_2624;
wire mux_o_2625;
wire mux_o_2626;
wire mux_o_2627;
wire mux_o_2628;
wire mux_o_2629;
wire mux_o_2630;
wire mux_o_2631;
wire mux_o_2632;
wire mux_o_2633;
wire mux_o_2634;
wire mux_o_2635;
wire mux_o_2636;
wire mux_o_2637;
wire mux_o_2638;
wire mux_o_2639;
wire mux_o_2640;
wire mux_o_2641;
wire mux_o_2642;
wire mux_o_2643;
wire mux_o_2644;
wire mux_o_2645;
wire mux_o_2646;
wire mux_o_2647;
wire mux_o_2648;
wire mux_o_2649;
wire mux_o_2650;
wire mux_o_2651;
wire mux_o_2652;
wire mux_o_2653;
wire mux_o_2654;
wire mux_o_2655;
wire mux_o_2656;
wire mux_o_2657;
wire mux_o_2658;
wire mux_o_2659;
wire mux_o_2660;
wire mux_o_2661;
wire mux_o_2662;
wire mux_o_2663;
wire mux_o_2664;
wire mux_o_2665;
wire mux_o_2667;
wire mux_o_2668;
wire mux_o_2669;
wire mux_o_2670;
wire mux_o_2671;
wire mux_o_2672;
wire mux_o_2673;
wire mux_o_2674;
wire mux_o_2675;
wire mux_o_2676;
wire mux_o_2677;
wire mux_o_2678;
wire mux_o_2679;
wire mux_o_2680;
wire mux_o_2681;
wire mux_o_2682;
wire mux_o_2683;
wire mux_o_2684;
wire mux_o_2685;
wire mux_o_2686;
wire mux_o_2687;
wire mux_o_2688;
wire mux_o_2689;
wire mux_o_2690;
wire mux_o_2691;
wire mux_o_2692;
wire mux_o_2693;
wire mux_o_2694;
wire mux_o_2695;
wire mux_o_2696;
wire mux_o_2697;
wire mux_o_2698;
wire mux_o_2699;
wire mux_o_2700;
wire mux_o_2701;
wire mux_o_2702;
wire mux_o_2703;
wire mux_o_2704;
wire mux_o_2705;
wire mux_o_2706;
wire mux_o_2707;
wire mux_o_2708;
wire mux_o_2709;
wire mux_o_2710;
wire mux_o_2711;
wire mux_o_2712;
wire mux_o_2713;
wire mux_o_2714;
wire mux_o_2715;
wire mux_o_2716;
wire mux_o_2717;
wire mux_o_2718;
wire mux_o_2719;
wire mux_o_2720;
wire mux_o_2721;
wire mux_o_2722;
wire mux_o_2723;
wire mux_o_2724;
wire mux_o_2725;
wire mux_o_2726;
wire mux_o_2727;
wire mux_o_2728;
wire mux_o_2729;
wire mux_o_2730;
wire mux_o_2731;
wire mux_o_2732;
wire mux_o_2733;
wire mux_o_2734;
wire mux_o_2735;
wire mux_o_2736;
wire mux_o_2737;
wire mux_o_2738;
wire mux_o_2739;
wire mux_o_2740;
wire mux_o_2741;
wire mux_o_2742;
wire mux_o_2743;
wire mux_o_2744;
wire mux_o_2745;
wire mux_o_2746;
wire mux_o_2747;
wire mux_o_2748;
wire mux_o_2749;
wire mux_o_2750;
wire mux_o_2751;
wire mux_o_2752;
wire mux_o_2753;
wire mux_o_2754;
wire mux_o_2755;
wire mux_o_2756;
wire mux_o_2757;
wire mux_o_2758;
wire mux_o_2759;
wire mux_o_2760;
wire mux_o_2761;
wire mux_o_2762;
wire mux_o_2763;
wire mux_o_2764;
wire mux_o_2765;
wire mux_o_2766;
wire mux_o_2767;
wire mux_o_2768;
wire mux_o_2769;
wire mux_o_2770;
wire mux_o_2771;
wire mux_o_2772;
wire mux_o_2773;
wire mux_o_2774;
wire mux_o_2775;
wire mux_o_2776;
wire mux_o_2777;
wire mux_o_2778;
wire mux_o_2779;
wire mux_o_2780;
wire mux_o_2781;
wire mux_o_2782;
wire mux_o_2783;
wire mux_o_2784;
wire mux_o_2785;
wire mux_o_2786;
wire mux_o_2787;
wire mux_o_2788;
wire mux_o_2789;
wire mux_o_2790;
wire mux_o_2791;
wire mux_o_2792;
wire mux_o_2794;
wire mux_o_2795;
wire mux_o_2796;
wire mux_o_2797;
wire mux_o_2798;
wire mux_o_2799;
wire mux_o_2800;
wire mux_o_2801;
wire mux_o_2802;
wire mux_o_2803;
wire mux_o_2804;
wire mux_o_2805;
wire mux_o_2806;
wire mux_o_2807;
wire mux_o_2808;
wire mux_o_2809;
wire mux_o_2810;
wire mux_o_2811;
wire mux_o_2812;
wire mux_o_2813;
wire mux_o_2814;
wire mux_o_2815;
wire mux_o_2816;
wire mux_o_2817;
wire mux_o_2818;
wire mux_o_2819;
wire mux_o_2820;
wire mux_o_2821;
wire mux_o_2822;
wire mux_o_2823;
wire mux_o_2824;
wire mux_o_2825;
wire mux_o_2826;
wire mux_o_2827;
wire mux_o_2828;
wire mux_o_2829;
wire mux_o_2830;
wire mux_o_2831;
wire mux_o_2832;
wire mux_o_2833;
wire mux_o_2834;
wire mux_o_2835;
wire mux_o_2836;
wire mux_o_2837;
wire mux_o_2838;
wire mux_o_2839;
wire mux_o_2840;
wire mux_o_2841;
wire mux_o_2842;
wire mux_o_2843;
wire mux_o_2844;
wire mux_o_2845;
wire mux_o_2846;
wire mux_o_2847;
wire mux_o_2848;
wire mux_o_2849;
wire mux_o_2850;
wire mux_o_2851;
wire mux_o_2852;
wire mux_o_2853;
wire mux_o_2854;
wire mux_o_2855;
wire mux_o_2856;
wire mux_o_2857;
wire mux_o_2858;
wire mux_o_2859;
wire mux_o_2860;
wire mux_o_2861;
wire mux_o_2862;
wire mux_o_2863;
wire mux_o_2864;
wire mux_o_2865;
wire mux_o_2866;
wire mux_o_2867;
wire mux_o_2868;
wire mux_o_2869;
wire mux_o_2870;
wire mux_o_2871;
wire mux_o_2872;
wire mux_o_2873;
wire mux_o_2874;
wire mux_o_2875;
wire mux_o_2876;
wire mux_o_2877;
wire mux_o_2878;
wire mux_o_2879;
wire mux_o_2880;
wire mux_o_2881;
wire mux_o_2882;
wire mux_o_2883;
wire mux_o_2884;
wire mux_o_2885;
wire mux_o_2886;
wire mux_o_2887;
wire mux_o_2888;
wire mux_o_2889;
wire mux_o_2890;
wire mux_o_2891;
wire mux_o_2892;
wire mux_o_2893;
wire mux_o_2894;
wire mux_o_2895;
wire mux_o_2896;
wire mux_o_2897;
wire mux_o_2898;
wire mux_o_2899;
wire mux_o_2900;
wire mux_o_2901;
wire mux_o_2902;
wire mux_o_2903;
wire mux_o_2904;
wire mux_o_2905;
wire mux_o_2906;
wire mux_o_2907;
wire mux_o_2908;
wire mux_o_2909;
wire mux_o_2910;
wire mux_o_2911;
wire mux_o_2912;
wire mux_o_2913;
wire mux_o_2914;
wire mux_o_2915;
wire mux_o_2916;
wire mux_o_2917;
wire mux_o_2918;
wire mux_o_2919;
wire mux_o_2921;
wire mux_o_2922;
wire mux_o_2923;
wire mux_o_2924;
wire mux_o_2925;
wire mux_o_2926;
wire mux_o_2927;
wire mux_o_2928;
wire mux_o_2929;
wire mux_o_2930;
wire mux_o_2931;
wire mux_o_2932;
wire mux_o_2933;
wire mux_o_2934;
wire mux_o_2935;
wire mux_o_2936;
wire mux_o_2937;
wire mux_o_2938;
wire mux_o_2939;
wire mux_o_2940;
wire mux_o_2941;
wire mux_o_2942;
wire mux_o_2943;
wire mux_o_2944;
wire mux_o_2945;
wire mux_o_2946;
wire mux_o_2947;
wire mux_o_2948;
wire mux_o_2949;
wire mux_o_2950;
wire mux_o_2951;
wire mux_o_2952;
wire mux_o_2953;
wire mux_o_2954;
wire mux_o_2955;
wire mux_o_2956;
wire mux_o_2957;
wire mux_o_2958;
wire mux_o_2959;
wire mux_o_2960;
wire mux_o_2961;
wire mux_o_2962;
wire mux_o_2963;
wire mux_o_2964;
wire mux_o_2965;
wire mux_o_2966;
wire mux_o_2967;
wire mux_o_2968;
wire mux_o_2969;
wire mux_o_2970;
wire mux_o_2971;
wire mux_o_2972;
wire mux_o_2973;
wire mux_o_2974;
wire mux_o_2975;
wire mux_o_2976;
wire mux_o_2977;
wire mux_o_2978;
wire mux_o_2979;
wire mux_o_2980;
wire mux_o_2981;
wire mux_o_2982;
wire mux_o_2983;
wire mux_o_2984;
wire mux_o_2985;
wire mux_o_2986;
wire mux_o_2987;
wire mux_o_2988;
wire mux_o_2989;
wire mux_o_2990;
wire mux_o_2991;
wire mux_o_2992;
wire mux_o_2993;
wire mux_o_2994;
wire mux_o_2995;
wire mux_o_2996;
wire mux_o_2997;
wire mux_o_2998;
wire mux_o_2999;
wire mux_o_3000;
wire mux_o_3001;
wire mux_o_3002;
wire mux_o_3003;
wire mux_o_3004;
wire mux_o_3005;
wire mux_o_3006;
wire mux_o_3007;
wire mux_o_3008;
wire mux_o_3009;
wire mux_o_3010;
wire mux_o_3011;
wire mux_o_3012;
wire mux_o_3013;
wire mux_o_3014;
wire mux_o_3015;
wire mux_o_3016;
wire mux_o_3017;
wire mux_o_3018;
wire mux_o_3019;
wire mux_o_3020;
wire mux_o_3021;
wire mux_o_3022;
wire mux_o_3023;
wire mux_o_3024;
wire mux_o_3025;
wire mux_o_3026;
wire mux_o_3027;
wire mux_o_3028;
wire mux_o_3029;
wire mux_o_3030;
wire mux_o_3031;
wire mux_o_3032;
wire mux_o_3033;
wire mux_o_3034;
wire mux_o_3035;
wire mux_o_3036;
wire mux_o_3037;
wire mux_o_3038;
wire mux_o_3039;
wire mux_o_3040;
wire mux_o_3041;
wire mux_o_3042;
wire mux_o_3043;
wire mux_o_3044;
wire mux_o_3045;
wire mux_o_3046;
wire mux_o_3048;
wire mux_o_3049;
wire mux_o_3050;
wire mux_o_3051;
wire mux_o_3052;
wire mux_o_3053;
wire mux_o_3054;
wire mux_o_3055;
wire mux_o_3056;
wire mux_o_3057;
wire mux_o_3058;
wire mux_o_3059;
wire mux_o_3060;
wire mux_o_3061;
wire mux_o_3062;
wire mux_o_3063;
wire mux_o_3064;
wire mux_o_3065;
wire mux_o_3066;
wire mux_o_3067;
wire mux_o_3068;
wire mux_o_3069;
wire mux_o_3070;
wire mux_o_3071;
wire mux_o_3072;
wire mux_o_3073;
wire mux_o_3074;
wire mux_o_3075;
wire mux_o_3076;
wire mux_o_3077;
wire mux_o_3078;
wire mux_o_3079;
wire mux_o_3080;
wire mux_o_3081;
wire mux_o_3082;
wire mux_o_3083;
wire mux_o_3084;
wire mux_o_3085;
wire mux_o_3086;
wire mux_o_3087;
wire mux_o_3088;
wire mux_o_3089;
wire mux_o_3090;
wire mux_o_3091;
wire mux_o_3092;
wire mux_o_3093;
wire mux_o_3094;
wire mux_o_3095;
wire mux_o_3096;
wire mux_o_3097;
wire mux_o_3098;
wire mux_o_3099;
wire mux_o_3100;
wire mux_o_3101;
wire mux_o_3102;
wire mux_o_3103;
wire mux_o_3104;
wire mux_o_3105;
wire mux_o_3106;
wire mux_o_3107;
wire mux_o_3108;
wire mux_o_3109;
wire mux_o_3110;
wire mux_o_3111;
wire mux_o_3112;
wire mux_o_3113;
wire mux_o_3114;
wire mux_o_3115;
wire mux_o_3116;
wire mux_o_3117;
wire mux_o_3118;
wire mux_o_3119;
wire mux_o_3120;
wire mux_o_3121;
wire mux_o_3122;
wire mux_o_3123;
wire mux_o_3124;
wire mux_o_3125;
wire mux_o_3126;
wire mux_o_3127;
wire mux_o_3128;
wire mux_o_3129;
wire mux_o_3130;
wire mux_o_3131;
wire mux_o_3132;
wire mux_o_3133;
wire mux_o_3134;
wire mux_o_3135;
wire mux_o_3136;
wire mux_o_3137;
wire mux_o_3138;
wire mux_o_3139;
wire mux_o_3140;
wire mux_o_3141;
wire mux_o_3142;
wire mux_o_3143;
wire mux_o_3144;
wire mux_o_3145;
wire mux_o_3146;
wire mux_o_3147;
wire mux_o_3148;
wire mux_o_3149;
wire mux_o_3150;
wire mux_o_3151;
wire mux_o_3152;
wire mux_o_3153;
wire mux_o_3154;
wire mux_o_3155;
wire mux_o_3156;
wire mux_o_3157;
wire mux_o_3158;
wire mux_o_3159;
wire mux_o_3160;
wire mux_o_3161;
wire mux_o_3162;
wire mux_o_3163;
wire mux_o_3164;
wire mux_o_3165;
wire mux_o_3166;
wire mux_o_3167;
wire mux_o_3168;
wire mux_o_3169;
wire mux_o_3170;
wire mux_o_3171;
wire mux_o_3172;
wire mux_o_3173;
wire mux_o_3175;
wire mux_o_3176;
wire mux_o_3177;
wire mux_o_3178;
wire mux_o_3179;
wire mux_o_3180;
wire mux_o_3181;
wire mux_o_3182;
wire mux_o_3183;
wire mux_o_3184;
wire mux_o_3185;
wire mux_o_3186;
wire mux_o_3187;
wire mux_o_3188;
wire mux_o_3189;
wire mux_o_3190;
wire mux_o_3191;
wire mux_o_3192;
wire mux_o_3193;
wire mux_o_3194;
wire mux_o_3195;
wire mux_o_3196;
wire mux_o_3197;
wire mux_o_3198;
wire mux_o_3199;
wire mux_o_3200;
wire mux_o_3201;
wire mux_o_3202;
wire mux_o_3203;
wire mux_o_3204;
wire mux_o_3205;
wire mux_o_3206;
wire mux_o_3207;
wire mux_o_3208;
wire mux_o_3209;
wire mux_o_3210;
wire mux_o_3211;
wire mux_o_3212;
wire mux_o_3213;
wire mux_o_3214;
wire mux_o_3215;
wire mux_o_3216;
wire mux_o_3217;
wire mux_o_3218;
wire mux_o_3219;
wire mux_o_3220;
wire mux_o_3221;
wire mux_o_3222;
wire mux_o_3223;
wire mux_o_3224;
wire mux_o_3225;
wire mux_o_3226;
wire mux_o_3227;
wire mux_o_3228;
wire mux_o_3229;
wire mux_o_3230;
wire mux_o_3231;
wire mux_o_3232;
wire mux_o_3233;
wire mux_o_3234;
wire mux_o_3235;
wire mux_o_3236;
wire mux_o_3237;
wire mux_o_3238;
wire mux_o_3239;
wire mux_o_3240;
wire mux_o_3241;
wire mux_o_3242;
wire mux_o_3243;
wire mux_o_3244;
wire mux_o_3245;
wire mux_o_3246;
wire mux_o_3247;
wire mux_o_3248;
wire mux_o_3249;
wire mux_o_3250;
wire mux_o_3251;
wire mux_o_3252;
wire mux_o_3253;
wire mux_o_3254;
wire mux_o_3255;
wire mux_o_3256;
wire mux_o_3257;
wire mux_o_3258;
wire mux_o_3259;
wire mux_o_3260;
wire mux_o_3261;
wire mux_o_3262;
wire mux_o_3263;
wire mux_o_3264;
wire mux_o_3265;
wire mux_o_3266;
wire mux_o_3267;
wire mux_o_3268;
wire mux_o_3269;
wire mux_o_3270;
wire mux_o_3271;
wire mux_o_3272;
wire mux_o_3273;
wire mux_o_3274;
wire mux_o_3275;
wire mux_o_3276;
wire mux_o_3277;
wire mux_o_3278;
wire mux_o_3279;
wire mux_o_3280;
wire mux_o_3281;
wire mux_o_3282;
wire mux_o_3283;
wire mux_o_3284;
wire mux_o_3285;
wire mux_o_3286;
wire mux_o_3287;
wire mux_o_3288;
wire mux_o_3289;
wire mux_o_3290;
wire mux_o_3291;
wire mux_o_3292;
wire mux_o_3293;
wire mux_o_3294;
wire mux_o_3295;
wire mux_o_3296;
wire mux_o_3297;
wire mux_o_3298;
wire mux_o_3299;
wire mux_o_3300;
wire mux_o_3302;
wire mux_o_3303;
wire mux_o_3304;
wire mux_o_3305;
wire mux_o_3306;
wire mux_o_3307;
wire mux_o_3308;
wire mux_o_3309;
wire mux_o_3310;
wire mux_o_3311;
wire mux_o_3312;
wire mux_o_3313;
wire mux_o_3314;
wire mux_o_3315;
wire mux_o_3316;
wire mux_o_3317;
wire mux_o_3318;
wire mux_o_3319;
wire mux_o_3320;
wire mux_o_3321;
wire mux_o_3322;
wire mux_o_3323;
wire mux_o_3324;
wire mux_o_3325;
wire mux_o_3326;
wire mux_o_3327;
wire mux_o_3328;
wire mux_o_3329;
wire mux_o_3330;
wire mux_o_3331;
wire mux_o_3332;
wire mux_o_3333;
wire mux_o_3334;
wire mux_o_3335;
wire mux_o_3336;
wire mux_o_3337;
wire mux_o_3338;
wire mux_o_3339;
wire mux_o_3340;
wire mux_o_3341;
wire mux_o_3342;
wire mux_o_3343;
wire mux_o_3344;
wire mux_o_3345;
wire mux_o_3346;
wire mux_o_3347;
wire mux_o_3348;
wire mux_o_3349;
wire mux_o_3350;
wire mux_o_3351;
wire mux_o_3352;
wire mux_o_3353;
wire mux_o_3354;
wire mux_o_3355;
wire mux_o_3356;
wire mux_o_3357;
wire mux_o_3358;
wire mux_o_3359;
wire mux_o_3360;
wire mux_o_3361;
wire mux_o_3362;
wire mux_o_3363;
wire mux_o_3364;
wire mux_o_3365;
wire mux_o_3366;
wire mux_o_3367;
wire mux_o_3368;
wire mux_o_3369;
wire mux_o_3370;
wire mux_o_3371;
wire mux_o_3372;
wire mux_o_3373;
wire mux_o_3374;
wire mux_o_3375;
wire mux_o_3376;
wire mux_o_3377;
wire mux_o_3378;
wire mux_o_3379;
wire mux_o_3380;
wire mux_o_3381;
wire mux_o_3382;
wire mux_o_3383;
wire mux_o_3384;
wire mux_o_3385;
wire mux_o_3386;
wire mux_o_3387;
wire mux_o_3388;
wire mux_o_3389;
wire mux_o_3390;
wire mux_o_3391;
wire mux_o_3392;
wire mux_o_3393;
wire mux_o_3394;
wire mux_o_3395;
wire mux_o_3396;
wire mux_o_3397;
wire mux_o_3398;
wire mux_o_3399;
wire mux_o_3400;
wire mux_o_3401;
wire mux_o_3402;
wire mux_o_3403;
wire mux_o_3404;
wire mux_o_3405;
wire mux_o_3406;
wire mux_o_3407;
wire mux_o_3408;
wire mux_o_3409;
wire mux_o_3410;
wire mux_o_3411;
wire mux_o_3412;
wire mux_o_3413;
wire mux_o_3414;
wire mux_o_3415;
wire mux_o_3416;
wire mux_o_3417;
wire mux_o_3418;
wire mux_o_3419;
wire mux_o_3420;
wire mux_o_3421;
wire mux_o_3422;
wire mux_o_3423;
wire mux_o_3424;
wire mux_o_3425;
wire mux_o_3426;
wire mux_o_3427;
wire mux_o_3429;
wire mux_o_3430;
wire mux_o_3431;
wire mux_o_3432;
wire mux_o_3433;
wire mux_o_3434;
wire mux_o_3435;
wire mux_o_3436;
wire mux_o_3437;
wire mux_o_3438;
wire mux_o_3439;
wire mux_o_3440;
wire mux_o_3441;
wire mux_o_3442;
wire mux_o_3443;
wire mux_o_3444;
wire mux_o_3445;
wire mux_o_3446;
wire mux_o_3447;
wire mux_o_3448;
wire mux_o_3449;
wire mux_o_3450;
wire mux_o_3451;
wire mux_o_3452;
wire mux_o_3453;
wire mux_o_3454;
wire mux_o_3455;
wire mux_o_3456;
wire mux_o_3457;
wire mux_o_3458;
wire mux_o_3459;
wire mux_o_3460;
wire mux_o_3461;
wire mux_o_3462;
wire mux_o_3463;
wire mux_o_3464;
wire mux_o_3465;
wire mux_o_3466;
wire mux_o_3467;
wire mux_o_3468;
wire mux_o_3469;
wire mux_o_3470;
wire mux_o_3471;
wire mux_o_3472;
wire mux_o_3473;
wire mux_o_3474;
wire mux_o_3475;
wire mux_o_3476;
wire mux_o_3477;
wire mux_o_3478;
wire mux_o_3479;
wire mux_o_3480;
wire mux_o_3481;
wire mux_o_3482;
wire mux_o_3483;
wire mux_o_3484;
wire mux_o_3485;
wire mux_o_3486;
wire mux_o_3487;
wire mux_o_3488;
wire mux_o_3489;
wire mux_o_3490;
wire mux_o_3491;
wire mux_o_3492;
wire mux_o_3493;
wire mux_o_3494;
wire mux_o_3495;
wire mux_o_3496;
wire mux_o_3497;
wire mux_o_3498;
wire mux_o_3499;
wire mux_o_3500;
wire mux_o_3501;
wire mux_o_3502;
wire mux_o_3503;
wire mux_o_3504;
wire mux_o_3505;
wire mux_o_3506;
wire mux_o_3507;
wire mux_o_3508;
wire mux_o_3509;
wire mux_o_3510;
wire mux_o_3511;
wire mux_o_3512;
wire mux_o_3513;
wire mux_o_3514;
wire mux_o_3515;
wire mux_o_3516;
wire mux_o_3517;
wire mux_o_3518;
wire mux_o_3519;
wire mux_o_3520;
wire mux_o_3521;
wire mux_o_3522;
wire mux_o_3523;
wire mux_o_3524;
wire mux_o_3525;
wire mux_o_3526;
wire mux_o_3527;
wire mux_o_3528;
wire mux_o_3529;
wire mux_o_3530;
wire mux_o_3531;
wire mux_o_3532;
wire mux_o_3533;
wire mux_o_3534;
wire mux_o_3535;
wire mux_o_3536;
wire mux_o_3537;
wire mux_o_3538;
wire mux_o_3539;
wire mux_o_3540;
wire mux_o_3541;
wire mux_o_3542;
wire mux_o_3543;
wire mux_o_3544;
wire mux_o_3545;
wire mux_o_3546;
wire mux_o_3547;
wire mux_o_3548;
wire mux_o_3549;
wire mux_o_3550;
wire mux_o_3551;
wire mux_o_3552;
wire mux_o_3553;
wire mux_o_3554;
wire mux_o_3556;
wire mux_o_3557;
wire mux_o_3558;
wire mux_o_3559;
wire mux_o_3560;
wire mux_o_3561;
wire mux_o_3562;
wire mux_o_3563;
wire mux_o_3564;
wire mux_o_3565;
wire mux_o_3566;
wire mux_o_3567;
wire mux_o_3568;
wire mux_o_3569;
wire mux_o_3570;
wire mux_o_3571;
wire mux_o_3572;
wire mux_o_3573;
wire mux_o_3574;
wire mux_o_3575;
wire mux_o_3576;
wire mux_o_3577;
wire mux_o_3578;
wire mux_o_3579;
wire mux_o_3580;
wire mux_o_3581;
wire mux_o_3582;
wire mux_o_3583;
wire mux_o_3584;
wire mux_o_3585;
wire mux_o_3586;
wire mux_o_3587;
wire mux_o_3588;
wire mux_o_3589;
wire mux_o_3590;
wire mux_o_3591;
wire mux_o_3592;
wire mux_o_3593;
wire mux_o_3594;
wire mux_o_3595;
wire mux_o_3596;
wire mux_o_3597;
wire mux_o_3598;
wire mux_o_3599;
wire mux_o_3600;
wire mux_o_3601;
wire mux_o_3602;
wire mux_o_3603;
wire mux_o_3604;
wire mux_o_3605;
wire mux_o_3606;
wire mux_o_3607;
wire mux_o_3608;
wire mux_o_3609;
wire mux_o_3610;
wire mux_o_3611;
wire mux_o_3612;
wire mux_o_3613;
wire mux_o_3614;
wire mux_o_3615;
wire mux_o_3616;
wire mux_o_3617;
wire mux_o_3618;
wire mux_o_3619;
wire mux_o_3620;
wire mux_o_3621;
wire mux_o_3622;
wire mux_o_3623;
wire mux_o_3624;
wire mux_o_3625;
wire mux_o_3626;
wire mux_o_3627;
wire mux_o_3628;
wire mux_o_3629;
wire mux_o_3630;
wire mux_o_3631;
wire mux_o_3632;
wire mux_o_3633;
wire mux_o_3634;
wire mux_o_3635;
wire mux_o_3636;
wire mux_o_3637;
wire mux_o_3638;
wire mux_o_3639;
wire mux_o_3640;
wire mux_o_3641;
wire mux_o_3642;
wire mux_o_3643;
wire mux_o_3644;
wire mux_o_3645;
wire mux_o_3646;
wire mux_o_3647;
wire mux_o_3648;
wire mux_o_3649;
wire mux_o_3650;
wire mux_o_3651;
wire mux_o_3652;
wire mux_o_3653;
wire mux_o_3654;
wire mux_o_3655;
wire mux_o_3656;
wire mux_o_3657;
wire mux_o_3658;
wire mux_o_3659;
wire mux_o_3660;
wire mux_o_3661;
wire mux_o_3662;
wire mux_o_3663;
wire mux_o_3664;
wire mux_o_3665;
wire mux_o_3666;
wire mux_o_3667;
wire mux_o_3668;
wire mux_o_3669;
wire mux_o_3670;
wire mux_o_3671;
wire mux_o_3672;
wire mux_o_3673;
wire mux_o_3674;
wire mux_o_3675;
wire mux_o_3676;
wire mux_o_3677;
wire mux_o_3678;
wire mux_o_3679;
wire mux_o_3680;
wire mux_o_3681;
wire mux_o_3683;
wire mux_o_3684;
wire mux_o_3685;
wire mux_o_3686;
wire mux_o_3687;
wire mux_o_3688;
wire mux_o_3689;
wire mux_o_3690;
wire mux_o_3691;
wire mux_o_3692;
wire mux_o_3693;
wire mux_o_3694;
wire mux_o_3695;
wire mux_o_3696;
wire mux_o_3697;
wire mux_o_3698;
wire mux_o_3699;
wire mux_o_3700;
wire mux_o_3701;
wire mux_o_3702;
wire mux_o_3703;
wire mux_o_3704;
wire mux_o_3705;
wire mux_o_3706;
wire mux_o_3707;
wire mux_o_3708;
wire mux_o_3709;
wire mux_o_3710;
wire mux_o_3711;
wire mux_o_3712;
wire mux_o_3713;
wire mux_o_3714;
wire mux_o_3715;
wire mux_o_3716;
wire mux_o_3717;
wire mux_o_3718;
wire mux_o_3719;
wire mux_o_3720;
wire mux_o_3721;
wire mux_o_3722;
wire mux_o_3723;
wire mux_o_3724;
wire mux_o_3725;
wire mux_o_3726;
wire mux_o_3727;
wire mux_o_3728;
wire mux_o_3729;
wire mux_o_3730;
wire mux_o_3731;
wire mux_o_3732;
wire mux_o_3733;
wire mux_o_3734;
wire mux_o_3735;
wire mux_o_3736;
wire mux_o_3737;
wire mux_o_3738;
wire mux_o_3739;
wire mux_o_3740;
wire mux_o_3741;
wire mux_o_3742;
wire mux_o_3743;
wire mux_o_3744;
wire mux_o_3745;
wire mux_o_3746;
wire mux_o_3747;
wire mux_o_3748;
wire mux_o_3749;
wire mux_o_3750;
wire mux_o_3751;
wire mux_o_3752;
wire mux_o_3753;
wire mux_o_3754;
wire mux_o_3755;
wire mux_o_3756;
wire mux_o_3757;
wire mux_o_3758;
wire mux_o_3759;
wire mux_o_3760;
wire mux_o_3761;
wire mux_o_3762;
wire mux_o_3763;
wire mux_o_3764;
wire mux_o_3765;
wire mux_o_3766;
wire mux_o_3767;
wire mux_o_3768;
wire mux_o_3769;
wire mux_o_3770;
wire mux_o_3771;
wire mux_o_3772;
wire mux_o_3773;
wire mux_o_3774;
wire mux_o_3775;
wire mux_o_3776;
wire mux_o_3777;
wire mux_o_3778;
wire mux_o_3779;
wire mux_o_3780;
wire mux_o_3781;
wire mux_o_3782;
wire mux_o_3783;
wire mux_o_3784;
wire mux_o_3785;
wire mux_o_3786;
wire mux_o_3787;
wire mux_o_3788;
wire mux_o_3789;
wire mux_o_3790;
wire mux_o_3791;
wire mux_o_3792;
wire mux_o_3793;
wire mux_o_3794;
wire mux_o_3795;
wire mux_o_3796;
wire mux_o_3797;
wire mux_o_3798;
wire mux_o_3799;
wire mux_o_3800;
wire mux_o_3801;
wire mux_o_3802;
wire mux_o_3803;
wire mux_o_3804;
wire mux_o_3805;
wire mux_o_3806;
wire mux_o_3807;
wire mux_o_3808;
wire mux_o_3810;
wire mux_o_3811;
wire mux_o_3812;
wire mux_o_3813;
wire mux_o_3814;
wire mux_o_3815;
wire mux_o_3816;
wire mux_o_3817;
wire mux_o_3818;
wire mux_o_3819;
wire mux_o_3820;
wire mux_o_3821;
wire mux_o_3822;
wire mux_o_3823;
wire mux_o_3824;
wire mux_o_3825;
wire mux_o_3826;
wire mux_o_3827;
wire mux_o_3828;
wire mux_o_3829;
wire mux_o_3830;
wire mux_o_3831;
wire mux_o_3832;
wire mux_o_3833;
wire mux_o_3834;
wire mux_o_3835;
wire mux_o_3836;
wire mux_o_3837;
wire mux_o_3838;
wire mux_o_3839;
wire mux_o_3840;
wire mux_o_3841;
wire mux_o_3842;
wire mux_o_3843;
wire mux_o_3844;
wire mux_o_3845;
wire mux_o_3846;
wire mux_o_3847;
wire mux_o_3848;
wire mux_o_3849;
wire mux_o_3850;
wire mux_o_3851;
wire mux_o_3852;
wire mux_o_3853;
wire mux_o_3854;
wire mux_o_3855;
wire mux_o_3856;
wire mux_o_3857;
wire mux_o_3858;
wire mux_o_3859;
wire mux_o_3860;
wire mux_o_3861;
wire mux_o_3862;
wire mux_o_3863;
wire mux_o_3864;
wire mux_o_3865;
wire mux_o_3866;
wire mux_o_3867;
wire mux_o_3868;
wire mux_o_3869;
wire mux_o_3870;
wire mux_o_3871;
wire mux_o_3872;
wire mux_o_3873;
wire mux_o_3874;
wire mux_o_3875;
wire mux_o_3876;
wire mux_o_3877;
wire mux_o_3878;
wire mux_o_3879;
wire mux_o_3880;
wire mux_o_3881;
wire mux_o_3882;
wire mux_o_3883;
wire mux_o_3884;
wire mux_o_3885;
wire mux_o_3886;
wire mux_o_3887;
wire mux_o_3888;
wire mux_o_3889;
wire mux_o_3890;
wire mux_o_3891;
wire mux_o_3892;
wire mux_o_3893;
wire mux_o_3894;
wire mux_o_3895;
wire mux_o_3896;
wire mux_o_3897;
wire mux_o_3898;
wire mux_o_3899;
wire mux_o_3900;
wire mux_o_3901;
wire mux_o_3902;
wire mux_o_3903;
wire mux_o_3904;
wire mux_o_3905;
wire mux_o_3906;
wire mux_o_3907;
wire mux_o_3908;
wire mux_o_3909;
wire mux_o_3910;
wire mux_o_3911;
wire mux_o_3912;
wire mux_o_3913;
wire mux_o_3914;
wire mux_o_3915;
wire mux_o_3916;
wire mux_o_3917;
wire mux_o_3918;
wire mux_o_3919;
wire mux_o_3920;
wire mux_o_3921;
wire mux_o_3922;
wire mux_o_3923;
wire mux_o_3924;
wire mux_o_3925;
wire mux_o_3926;
wire mux_o_3927;
wire mux_o_3928;
wire mux_o_3929;
wire mux_o_3930;
wire mux_o_3931;
wire mux_o_3932;
wire mux_o_3933;
wire mux_o_3934;
wire mux_o_3935;
wire mux_o_3937;
wire mux_o_3938;
wire mux_o_3939;
wire mux_o_3940;
wire mux_o_3941;
wire mux_o_3942;
wire mux_o_3943;
wire mux_o_3944;
wire mux_o_3945;
wire mux_o_3946;
wire mux_o_3947;
wire mux_o_3948;
wire mux_o_3949;
wire mux_o_3950;
wire mux_o_3951;
wire mux_o_3952;
wire mux_o_3953;
wire mux_o_3954;
wire mux_o_3955;
wire mux_o_3956;
wire mux_o_3957;
wire mux_o_3958;
wire mux_o_3959;
wire mux_o_3960;
wire mux_o_3961;
wire mux_o_3962;
wire mux_o_3963;
wire mux_o_3964;
wire mux_o_3965;
wire mux_o_3966;
wire mux_o_3967;
wire mux_o_3968;
wire mux_o_3969;
wire mux_o_3970;
wire mux_o_3971;
wire mux_o_3972;
wire mux_o_3973;
wire mux_o_3974;
wire mux_o_3975;
wire mux_o_3976;
wire mux_o_3977;
wire mux_o_3978;
wire mux_o_3979;
wire mux_o_3980;
wire mux_o_3981;
wire mux_o_3982;
wire mux_o_3983;
wire mux_o_3984;
wire mux_o_3985;
wire mux_o_3986;
wire mux_o_3987;
wire mux_o_3988;
wire mux_o_3989;
wire mux_o_3990;
wire mux_o_3991;
wire mux_o_3992;
wire mux_o_3993;
wire mux_o_3994;
wire mux_o_3995;
wire mux_o_3996;
wire mux_o_3997;
wire mux_o_3998;
wire mux_o_3999;
wire mux_o_4000;
wire mux_o_4001;
wire mux_o_4002;
wire mux_o_4003;
wire mux_o_4004;
wire mux_o_4005;
wire mux_o_4006;
wire mux_o_4007;
wire mux_o_4008;
wire mux_o_4009;
wire mux_o_4010;
wire mux_o_4011;
wire mux_o_4012;
wire mux_o_4013;
wire mux_o_4014;
wire mux_o_4015;
wire mux_o_4016;
wire mux_o_4017;
wire mux_o_4018;
wire mux_o_4019;
wire mux_o_4020;
wire mux_o_4021;
wire mux_o_4022;
wire mux_o_4023;
wire mux_o_4024;
wire mux_o_4025;
wire mux_o_4026;
wire mux_o_4027;
wire mux_o_4028;
wire mux_o_4029;
wire mux_o_4030;
wire mux_o_4031;
wire mux_o_4032;
wire mux_o_4033;
wire mux_o_4034;
wire mux_o_4035;
wire mux_o_4036;
wire mux_o_4037;
wire mux_o_4038;
wire mux_o_4039;
wire mux_o_4040;
wire mux_o_4041;
wire mux_o_4042;
wire mux_o_4043;
wire mux_o_4044;
wire mux_o_4045;
wire mux_o_4046;
wire mux_o_4047;
wire mux_o_4048;
wire mux_o_4049;
wire mux_o_4050;
wire mux_o_4051;
wire mux_o_4052;
wire mux_o_4053;
wire mux_o_4054;
wire mux_o_4055;
wire mux_o_4056;
wire mux_o_4057;
wire mux_o_4058;
wire mux_o_4059;
wire mux_o_4060;
wire mux_o_4061;
wire mux_o_4062;
wire gw_vcc;

assign gw_vcc = 1'b1;

INV inv_inst_0 (.I(wad[4]), .O(wad4_inv));

INV inv_inst_1 (.I(wad[5]), .O(wad5_inv));

INV inv_inst_2 (.I(wad[6]), .O(wad6_inv));

INV inv_inst_3 (.I(wad[7]), .O(wad7_inv));

INV inv_inst_4 (.I(wad[8]), .O(wad8_inv));

INV inv_inst_5 (.I(wad[9]), .O(wad9_inv));

INV inv_inst_6 (.I(wad[10]), .O(wad10_inv));

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_0.INIT = 16'h8000;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_1.INIT = 16'h8000;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(lut_f_0),
  .I1(lut_f_1),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_2.INIT = 16'h8000;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_3.INIT = 16'h8000;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_4.INIT = 16'h8000;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(lut_f_3),
  .I1(lut_f_4),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_5.INIT = 16'h8000;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_6.INIT = 16'h8000;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_7.INIT = 16'h8000;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(lut_f_6),
  .I1(lut_f_7),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_8.INIT = 16'h8000;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_9.INIT = 16'h8000;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_10.INIT = 16'h8000;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(lut_f_9),
  .I1(lut_f_10),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_11.INIT = 16'h8000;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_12.INIT = 16'h8000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_13.INIT = 16'h8000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(lut_f_12),
  .I1(lut_f_13),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_14.INIT = 16'h8000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_15.INIT = 16'h8000;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_16.INIT = 16'h8000;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(lut_f_15),
  .I1(lut_f_16),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_17.INIT = 16'h8000;
LUT4 lut_inst_18 (
  .F(lut_f_18),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_18.INIT = 16'h8000;
LUT4 lut_inst_19 (
  .F(lut_f_19),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_19.INIT = 16'h8000;
LUT4 lut_inst_20 (
  .F(lut_f_20),
  .I0(lut_f_18),
  .I1(lut_f_19),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_20.INIT = 16'h8000;
LUT4 lut_inst_21 (
  .F(lut_f_21),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_21.INIT = 16'h8000;
LUT4 lut_inst_22 (
  .F(lut_f_22),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_22.INIT = 16'h8000;
LUT4 lut_inst_23 (
  .F(lut_f_23),
  .I0(lut_f_21),
  .I1(lut_f_22),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_23.INIT = 16'h8000;
LUT4 lut_inst_24 (
  .F(lut_f_24),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_24.INIT = 16'h8000;
LUT4 lut_inst_25 (
  .F(lut_f_25),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_25.INIT = 16'h8000;
LUT4 lut_inst_26 (
  .F(lut_f_26),
  .I0(lut_f_24),
  .I1(lut_f_25),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_26.INIT = 16'h8000;
LUT4 lut_inst_27 (
  .F(lut_f_27),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_27.INIT = 16'h8000;
LUT4 lut_inst_28 (
  .F(lut_f_28),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_28.INIT = 16'h8000;
LUT4 lut_inst_29 (
  .F(lut_f_29),
  .I0(lut_f_27),
  .I1(lut_f_28),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_29.INIT = 16'h8000;
LUT4 lut_inst_30 (
  .F(lut_f_30),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_30.INIT = 16'h8000;
LUT4 lut_inst_31 (
  .F(lut_f_31),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_31.INIT = 16'h8000;
LUT4 lut_inst_32 (
  .F(lut_f_32),
  .I0(lut_f_30),
  .I1(lut_f_31),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_32.INIT = 16'h8000;
LUT4 lut_inst_33 (
  .F(lut_f_33),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_33.INIT = 16'h8000;
LUT4 lut_inst_34 (
  .F(lut_f_34),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_34.INIT = 16'h8000;
LUT4 lut_inst_35 (
  .F(lut_f_35),
  .I0(lut_f_33),
  .I1(lut_f_34),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_35.INIT = 16'h8000;
LUT4 lut_inst_36 (
  .F(lut_f_36),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_36.INIT = 16'h8000;
LUT4 lut_inst_37 (
  .F(lut_f_37),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_37.INIT = 16'h8000;
LUT4 lut_inst_38 (
  .F(lut_f_38),
  .I0(lut_f_36),
  .I1(lut_f_37),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_38.INIT = 16'h8000;
LUT4 lut_inst_39 (
  .F(lut_f_39),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_39.INIT = 16'h8000;
LUT4 lut_inst_40 (
  .F(lut_f_40),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_40.INIT = 16'h8000;
LUT4 lut_inst_41 (
  .F(lut_f_41),
  .I0(lut_f_39),
  .I1(lut_f_40),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_41.INIT = 16'h8000;
LUT4 lut_inst_42 (
  .F(lut_f_42),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_42.INIT = 16'h8000;
LUT4 lut_inst_43 (
  .F(lut_f_43),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_43.INIT = 16'h8000;
LUT4 lut_inst_44 (
  .F(lut_f_44),
  .I0(lut_f_42),
  .I1(lut_f_43),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_44.INIT = 16'h8000;
LUT4 lut_inst_45 (
  .F(lut_f_45),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_45.INIT = 16'h8000;
LUT4 lut_inst_46 (
  .F(lut_f_46),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_46.INIT = 16'h8000;
LUT4 lut_inst_47 (
  .F(lut_f_47),
  .I0(lut_f_45),
  .I1(lut_f_46),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_47.INIT = 16'h8000;
LUT4 lut_inst_48 (
  .F(lut_f_48),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_48.INIT = 16'h8000;
LUT4 lut_inst_49 (
  .F(lut_f_49),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_49.INIT = 16'h8000;
LUT4 lut_inst_50 (
  .F(lut_f_50),
  .I0(lut_f_48),
  .I1(lut_f_49),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_50.INIT = 16'h8000;
LUT4 lut_inst_51 (
  .F(lut_f_51),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_51.INIT = 16'h8000;
LUT4 lut_inst_52 (
  .F(lut_f_52),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_52.INIT = 16'h8000;
LUT4 lut_inst_53 (
  .F(lut_f_53),
  .I0(lut_f_51),
  .I1(lut_f_52),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_53.INIT = 16'h8000;
LUT4 lut_inst_54 (
  .F(lut_f_54),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_54.INIT = 16'h8000;
LUT4 lut_inst_55 (
  .F(lut_f_55),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_55.INIT = 16'h8000;
LUT4 lut_inst_56 (
  .F(lut_f_56),
  .I0(lut_f_54),
  .I1(lut_f_55),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_56.INIT = 16'h8000;
LUT4 lut_inst_57 (
  .F(lut_f_57),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_57.INIT = 16'h8000;
LUT4 lut_inst_58 (
  .F(lut_f_58),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_58.INIT = 16'h8000;
LUT4 lut_inst_59 (
  .F(lut_f_59),
  .I0(lut_f_57),
  .I1(lut_f_58),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_59.INIT = 16'h8000;
LUT4 lut_inst_60 (
  .F(lut_f_60),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_60.INIT = 16'h8000;
LUT4 lut_inst_61 (
  .F(lut_f_61),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_61.INIT = 16'h8000;
LUT4 lut_inst_62 (
  .F(lut_f_62),
  .I0(lut_f_60),
  .I1(lut_f_61),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_62.INIT = 16'h8000;
LUT4 lut_inst_63 (
  .F(lut_f_63),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_63.INIT = 16'h8000;
LUT4 lut_inst_64 (
  .F(lut_f_64),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_64.INIT = 16'h8000;
LUT4 lut_inst_65 (
  .F(lut_f_65),
  .I0(lut_f_63),
  .I1(lut_f_64),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_65.INIT = 16'h8000;
LUT4 lut_inst_66 (
  .F(lut_f_66),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_66.INIT = 16'h8000;
LUT4 lut_inst_67 (
  .F(lut_f_67),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_67.INIT = 16'h8000;
LUT4 lut_inst_68 (
  .F(lut_f_68),
  .I0(lut_f_66),
  .I1(lut_f_67),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_68.INIT = 16'h8000;
LUT4 lut_inst_69 (
  .F(lut_f_69),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_69.INIT = 16'h8000;
LUT4 lut_inst_70 (
  .F(lut_f_70),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_70.INIT = 16'h8000;
LUT4 lut_inst_71 (
  .F(lut_f_71),
  .I0(lut_f_69),
  .I1(lut_f_70),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_71.INIT = 16'h8000;
LUT4 lut_inst_72 (
  .F(lut_f_72),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_72.INIT = 16'h8000;
LUT4 lut_inst_73 (
  .F(lut_f_73),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_73.INIT = 16'h8000;
LUT4 lut_inst_74 (
  .F(lut_f_74),
  .I0(lut_f_72),
  .I1(lut_f_73),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_74.INIT = 16'h8000;
LUT4 lut_inst_75 (
  .F(lut_f_75),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_75.INIT = 16'h8000;
LUT4 lut_inst_76 (
  .F(lut_f_76),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_76.INIT = 16'h8000;
LUT4 lut_inst_77 (
  .F(lut_f_77),
  .I0(lut_f_75),
  .I1(lut_f_76),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_77.INIT = 16'h8000;
LUT4 lut_inst_78 (
  .F(lut_f_78),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_78.INIT = 16'h8000;
LUT4 lut_inst_79 (
  .F(lut_f_79),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_79.INIT = 16'h8000;
LUT4 lut_inst_80 (
  .F(lut_f_80),
  .I0(lut_f_78),
  .I1(lut_f_79),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_80.INIT = 16'h8000;
LUT4 lut_inst_81 (
  .F(lut_f_81),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_81.INIT = 16'h8000;
LUT4 lut_inst_82 (
  .F(lut_f_82),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_82.INIT = 16'h8000;
LUT4 lut_inst_83 (
  .F(lut_f_83),
  .I0(lut_f_81),
  .I1(lut_f_82),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_83.INIT = 16'h8000;
LUT4 lut_inst_84 (
  .F(lut_f_84),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_84.INIT = 16'h8000;
LUT4 lut_inst_85 (
  .F(lut_f_85),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_85.INIT = 16'h8000;
LUT4 lut_inst_86 (
  .F(lut_f_86),
  .I0(lut_f_84),
  .I1(lut_f_85),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_86.INIT = 16'h8000;
LUT4 lut_inst_87 (
  .F(lut_f_87),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_87.INIT = 16'h8000;
LUT4 lut_inst_88 (
  .F(lut_f_88),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_88.INIT = 16'h8000;
LUT4 lut_inst_89 (
  .F(lut_f_89),
  .I0(lut_f_87),
  .I1(lut_f_88),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_89.INIT = 16'h8000;
LUT4 lut_inst_90 (
  .F(lut_f_90),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_90.INIT = 16'h8000;
LUT4 lut_inst_91 (
  .F(lut_f_91),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_91.INIT = 16'h8000;
LUT4 lut_inst_92 (
  .F(lut_f_92),
  .I0(lut_f_90),
  .I1(lut_f_91),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_92.INIT = 16'h8000;
LUT4 lut_inst_93 (
  .F(lut_f_93),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_93.INIT = 16'h8000;
LUT4 lut_inst_94 (
  .F(lut_f_94),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad10_inv)
);
defparam lut_inst_94.INIT = 16'h8000;
LUT4 lut_inst_95 (
  .F(lut_f_95),
  .I0(lut_f_93),
  .I1(lut_f_94),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_95.INIT = 16'h8000;
LUT4 lut_inst_96 (
  .F(lut_f_96),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_96.INIT = 16'h8000;
LUT4 lut_inst_97 (
  .F(lut_f_97),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_97.INIT = 16'h8000;
LUT4 lut_inst_98 (
  .F(lut_f_98),
  .I0(lut_f_96),
  .I1(lut_f_97),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_98.INIT = 16'h8000;
LUT4 lut_inst_99 (
  .F(lut_f_99),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_99.INIT = 16'h8000;
LUT4 lut_inst_100 (
  .F(lut_f_100),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_100.INIT = 16'h8000;
LUT4 lut_inst_101 (
  .F(lut_f_101),
  .I0(lut_f_99),
  .I1(lut_f_100),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_101.INIT = 16'h8000;
LUT4 lut_inst_102 (
  .F(lut_f_102),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_102.INIT = 16'h8000;
LUT4 lut_inst_103 (
  .F(lut_f_103),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_103.INIT = 16'h8000;
LUT4 lut_inst_104 (
  .F(lut_f_104),
  .I0(lut_f_102),
  .I1(lut_f_103),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_104.INIT = 16'h8000;
LUT4 lut_inst_105 (
  .F(lut_f_105),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_105.INIT = 16'h8000;
LUT4 lut_inst_106 (
  .F(lut_f_106),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_106.INIT = 16'h8000;
LUT4 lut_inst_107 (
  .F(lut_f_107),
  .I0(lut_f_105),
  .I1(lut_f_106),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_107.INIT = 16'h8000;
LUT4 lut_inst_108 (
  .F(lut_f_108),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_108.INIT = 16'h8000;
LUT4 lut_inst_109 (
  .F(lut_f_109),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_109.INIT = 16'h8000;
LUT4 lut_inst_110 (
  .F(lut_f_110),
  .I0(lut_f_108),
  .I1(lut_f_109),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_110.INIT = 16'h8000;
LUT4 lut_inst_111 (
  .F(lut_f_111),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_111.INIT = 16'h8000;
LUT4 lut_inst_112 (
  .F(lut_f_112),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_112.INIT = 16'h8000;
LUT4 lut_inst_113 (
  .F(lut_f_113),
  .I0(lut_f_111),
  .I1(lut_f_112),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_113.INIT = 16'h8000;
LUT4 lut_inst_114 (
  .F(lut_f_114),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_114.INIT = 16'h8000;
LUT4 lut_inst_115 (
  .F(lut_f_115),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_115.INIT = 16'h8000;
LUT4 lut_inst_116 (
  .F(lut_f_116),
  .I0(lut_f_114),
  .I1(lut_f_115),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_116.INIT = 16'h8000;
LUT4 lut_inst_117 (
  .F(lut_f_117),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_117.INIT = 16'h8000;
LUT4 lut_inst_118 (
  .F(lut_f_118),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_118.INIT = 16'h8000;
LUT4 lut_inst_119 (
  .F(lut_f_119),
  .I0(lut_f_117),
  .I1(lut_f_118),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_119.INIT = 16'h8000;
LUT4 lut_inst_120 (
  .F(lut_f_120),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_120.INIT = 16'h8000;
LUT4 lut_inst_121 (
  .F(lut_f_121),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_121.INIT = 16'h8000;
LUT4 lut_inst_122 (
  .F(lut_f_122),
  .I0(lut_f_120),
  .I1(lut_f_121),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_122.INIT = 16'h8000;
LUT4 lut_inst_123 (
  .F(lut_f_123),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_123.INIT = 16'h8000;
LUT4 lut_inst_124 (
  .F(lut_f_124),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_124.INIT = 16'h8000;
LUT4 lut_inst_125 (
  .F(lut_f_125),
  .I0(lut_f_123),
  .I1(lut_f_124),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_125.INIT = 16'h8000;
LUT4 lut_inst_126 (
  .F(lut_f_126),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_126.INIT = 16'h8000;
LUT4 lut_inst_127 (
  .F(lut_f_127),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_127.INIT = 16'h8000;
LUT4 lut_inst_128 (
  .F(lut_f_128),
  .I0(lut_f_126),
  .I1(lut_f_127),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_128.INIT = 16'h8000;
LUT4 lut_inst_129 (
  .F(lut_f_129),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_129.INIT = 16'h8000;
LUT4 lut_inst_130 (
  .F(lut_f_130),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_130.INIT = 16'h8000;
LUT4 lut_inst_131 (
  .F(lut_f_131),
  .I0(lut_f_129),
  .I1(lut_f_130),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_131.INIT = 16'h8000;
LUT4 lut_inst_132 (
  .F(lut_f_132),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_132.INIT = 16'h8000;
LUT4 lut_inst_133 (
  .F(lut_f_133),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_133.INIT = 16'h8000;
LUT4 lut_inst_134 (
  .F(lut_f_134),
  .I0(lut_f_132),
  .I1(lut_f_133),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_134.INIT = 16'h8000;
LUT4 lut_inst_135 (
  .F(lut_f_135),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_135.INIT = 16'h8000;
LUT4 lut_inst_136 (
  .F(lut_f_136),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_136.INIT = 16'h8000;
LUT4 lut_inst_137 (
  .F(lut_f_137),
  .I0(lut_f_135),
  .I1(lut_f_136),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_137.INIT = 16'h8000;
LUT4 lut_inst_138 (
  .F(lut_f_138),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_138.INIT = 16'h8000;
LUT4 lut_inst_139 (
  .F(lut_f_139),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_139.INIT = 16'h8000;
LUT4 lut_inst_140 (
  .F(lut_f_140),
  .I0(lut_f_138),
  .I1(lut_f_139),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_140.INIT = 16'h8000;
LUT4 lut_inst_141 (
  .F(lut_f_141),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_141.INIT = 16'h8000;
LUT4 lut_inst_142 (
  .F(lut_f_142),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_142.INIT = 16'h8000;
LUT4 lut_inst_143 (
  .F(lut_f_143),
  .I0(lut_f_141),
  .I1(lut_f_142),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_143.INIT = 16'h8000;
LUT4 lut_inst_144 (
  .F(lut_f_144),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_144.INIT = 16'h8000;
LUT4 lut_inst_145 (
  .F(lut_f_145),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_145.INIT = 16'h8000;
LUT4 lut_inst_146 (
  .F(lut_f_146),
  .I0(lut_f_144),
  .I1(lut_f_145),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_146.INIT = 16'h8000;
LUT4 lut_inst_147 (
  .F(lut_f_147),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_147.INIT = 16'h8000;
LUT4 lut_inst_148 (
  .F(lut_f_148),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_148.INIT = 16'h8000;
LUT4 lut_inst_149 (
  .F(lut_f_149),
  .I0(lut_f_147),
  .I1(lut_f_148),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_149.INIT = 16'h8000;
LUT4 lut_inst_150 (
  .F(lut_f_150),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_150.INIT = 16'h8000;
LUT4 lut_inst_151 (
  .F(lut_f_151),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_151.INIT = 16'h8000;
LUT4 lut_inst_152 (
  .F(lut_f_152),
  .I0(lut_f_150),
  .I1(lut_f_151),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_152.INIT = 16'h8000;
LUT4 lut_inst_153 (
  .F(lut_f_153),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_153.INIT = 16'h8000;
LUT4 lut_inst_154 (
  .F(lut_f_154),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_154.INIT = 16'h8000;
LUT4 lut_inst_155 (
  .F(lut_f_155),
  .I0(lut_f_153),
  .I1(lut_f_154),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_155.INIT = 16'h8000;
LUT4 lut_inst_156 (
  .F(lut_f_156),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_156.INIT = 16'h8000;
LUT4 lut_inst_157 (
  .F(lut_f_157),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_157.INIT = 16'h8000;
LUT4 lut_inst_158 (
  .F(lut_f_158),
  .I0(lut_f_156),
  .I1(lut_f_157),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_158.INIT = 16'h8000;
LUT4 lut_inst_159 (
  .F(lut_f_159),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_159.INIT = 16'h8000;
LUT4 lut_inst_160 (
  .F(lut_f_160),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_160.INIT = 16'h8000;
LUT4 lut_inst_161 (
  .F(lut_f_161),
  .I0(lut_f_159),
  .I1(lut_f_160),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_161.INIT = 16'h8000;
LUT4 lut_inst_162 (
  .F(lut_f_162),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_162.INIT = 16'h8000;
LUT4 lut_inst_163 (
  .F(lut_f_163),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_163.INIT = 16'h8000;
LUT4 lut_inst_164 (
  .F(lut_f_164),
  .I0(lut_f_162),
  .I1(lut_f_163),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_164.INIT = 16'h8000;
LUT4 lut_inst_165 (
  .F(lut_f_165),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_165.INIT = 16'h8000;
LUT4 lut_inst_166 (
  .F(lut_f_166),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_166.INIT = 16'h8000;
LUT4 lut_inst_167 (
  .F(lut_f_167),
  .I0(lut_f_165),
  .I1(lut_f_166),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_167.INIT = 16'h8000;
LUT4 lut_inst_168 (
  .F(lut_f_168),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_168.INIT = 16'h8000;
LUT4 lut_inst_169 (
  .F(lut_f_169),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_169.INIT = 16'h8000;
LUT4 lut_inst_170 (
  .F(lut_f_170),
  .I0(lut_f_168),
  .I1(lut_f_169),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_170.INIT = 16'h8000;
LUT4 lut_inst_171 (
  .F(lut_f_171),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_171.INIT = 16'h8000;
LUT4 lut_inst_172 (
  .F(lut_f_172),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_172.INIT = 16'h8000;
LUT4 lut_inst_173 (
  .F(lut_f_173),
  .I0(lut_f_171),
  .I1(lut_f_172),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_173.INIT = 16'h8000;
LUT4 lut_inst_174 (
  .F(lut_f_174),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_174.INIT = 16'h8000;
LUT4 lut_inst_175 (
  .F(lut_f_175),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_175.INIT = 16'h8000;
LUT4 lut_inst_176 (
  .F(lut_f_176),
  .I0(lut_f_174),
  .I1(lut_f_175),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_176.INIT = 16'h8000;
LUT4 lut_inst_177 (
  .F(lut_f_177),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_177.INIT = 16'h8000;
LUT4 lut_inst_178 (
  .F(lut_f_178),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_178.INIT = 16'h8000;
LUT4 lut_inst_179 (
  .F(lut_f_179),
  .I0(lut_f_177),
  .I1(lut_f_178),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_179.INIT = 16'h8000;
LUT4 lut_inst_180 (
  .F(lut_f_180),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_180.INIT = 16'h8000;
LUT4 lut_inst_181 (
  .F(lut_f_181),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_181.INIT = 16'h8000;
LUT4 lut_inst_182 (
  .F(lut_f_182),
  .I0(lut_f_180),
  .I1(lut_f_181),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_182.INIT = 16'h8000;
LUT4 lut_inst_183 (
  .F(lut_f_183),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_183.INIT = 16'h8000;
LUT4 lut_inst_184 (
  .F(lut_f_184),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_184.INIT = 16'h8000;
LUT4 lut_inst_185 (
  .F(lut_f_185),
  .I0(lut_f_183),
  .I1(lut_f_184),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_185.INIT = 16'h8000;
LUT4 lut_inst_186 (
  .F(lut_f_186),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_186.INIT = 16'h8000;
LUT4 lut_inst_187 (
  .F(lut_f_187),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_187.INIT = 16'h8000;
LUT4 lut_inst_188 (
  .F(lut_f_188),
  .I0(lut_f_186),
  .I1(lut_f_187),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_188.INIT = 16'h8000;
LUT4 lut_inst_189 (
  .F(lut_f_189),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_189.INIT = 16'h8000;
LUT4 lut_inst_190 (
  .F(lut_f_190),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad10_inv)
);
defparam lut_inst_190.INIT = 16'h8000;
LUT4 lut_inst_191 (
  .F(lut_f_191),
  .I0(lut_f_189),
  .I1(lut_f_190),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_191.INIT = 16'h8000;
LUT4 lut_inst_192 (
  .F(lut_f_192),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_192.INIT = 16'h8000;
LUT4 lut_inst_193 (
  .F(lut_f_193),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_193.INIT = 16'h8000;
LUT4 lut_inst_194 (
  .F(lut_f_194),
  .I0(lut_f_192),
  .I1(lut_f_193),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_194.INIT = 16'h8000;
LUT4 lut_inst_195 (
  .F(lut_f_195),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_195.INIT = 16'h8000;
LUT4 lut_inst_196 (
  .F(lut_f_196),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_196.INIT = 16'h8000;
LUT4 lut_inst_197 (
  .F(lut_f_197),
  .I0(lut_f_195),
  .I1(lut_f_196),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_197.INIT = 16'h8000;
LUT4 lut_inst_198 (
  .F(lut_f_198),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_198.INIT = 16'h8000;
LUT4 lut_inst_199 (
  .F(lut_f_199),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_199.INIT = 16'h8000;
LUT4 lut_inst_200 (
  .F(lut_f_200),
  .I0(lut_f_198),
  .I1(lut_f_199),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_200.INIT = 16'h8000;
LUT4 lut_inst_201 (
  .F(lut_f_201),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_201.INIT = 16'h8000;
LUT4 lut_inst_202 (
  .F(lut_f_202),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_202.INIT = 16'h8000;
LUT4 lut_inst_203 (
  .F(lut_f_203),
  .I0(lut_f_201),
  .I1(lut_f_202),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_203.INIT = 16'h8000;
LUT4 lut_inst_204 (
  .F(lut_f_204),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_204.INIT = 16'h8000;
LUT4 lut_inst_205 (
  .F(lut_f_205),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_205.INIT = 16'h8000;
LUT4 lut_inst_206 (
  .F(lut_f_206),
  .I0(lut_f_204),
  .I1(lut_f_205),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_206.INIT = 16'h8000;
LUT4 lut_inst_207 (
  .F(lut_f_207),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_207.INIT = 16'h8000;
LUT4 lut_inst_208 (
  .F(lut_f_208),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_208.INIT = 16'h8000;
LUT4 lut_inst_209 (
  .F(lut_f_209),
  .I0(lut_f_207),
  .I1(lut_f_208),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_209.INIT = 16'h8000;
LUT4 lut_inst_210 (
  .F(lut_f_210),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_210.INIT = 16'h8000;
LUT4 lut_inst_211 (
  .F(lut_f_211),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_211.INIT = 16'h8000;
LUT4 lut_inst_212 (
  .F(lut_f_212),
  .I0(lut_f_210),
  .I1(lut_f_211),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_212.INIT = 16'h8000;
LUT4 lut_inst_213 (
  .F(lut_f_213),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_213.INIT = 16'h8000;
LUT4 lut_inst_214 (
  .F(lut_f_214),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_214.INIT = 16'h8000;
LUT4 lut_inst_215 (
  .F(lut_f_215),
  .I0(lut_f_213),
  .I1(lut_f_214),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_215.INIT = 16'h8000;
LUT4 lut_inst_216 (
  .F(lut_f_216),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_216.INIT = 16'h8000;
LUT4 lut_inst_217 (
  .F(lut_f_217),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_217.INIT = 16'h8000;
LUT4 lut_inst_218 (
  .F(lut_f_218),
  .I0(lut_f_216),
  .I1(lut_f_217),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_218.INIT = 16'h8000;
LUT4 lut_inst_219 (
  .F(lut_f_219),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_219.INIT = 16'h8000;
LUT4 lut_inst_220 (
  .F(lut_f_220),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_220.INIT = 16'h8000;
LUT4 lut_inst_221 (
  .F(lut_f_221),
  .I0(lut_f_219),
  .I1(lut_f_220),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_221.INIT = 16'h8000;
LUT4 lut_inst_222 (
  .F(lut_f_222),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_222.INIT = 16'h8000;
LUT4 lut_inst_223 (
  .F(lut_f_223),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_223.INIT = 16'h8000;
LUT4 lut_inst_224 (
  .F(lut_f_224),
  .I0(lut_f_222),
  .I1(lut_f_223),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_224.INIT = 16'h8000;
LUT4 lut_inst_225 (
  .F(lut_f_225),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_225.INIT = 16'h8000;
LUT4 lut_inst_226 (
  .F(lut_f_226),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_226.INIT = 16'h8000;
LUT4 lut_inst_227 (
  .F(lut_f_227),
  .I0(lut_f_225),
  .I1(lut_f_226),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_227.INIT = 16'h8000;
LUT4 lut_inst_228 (
  .F(lut_f_228),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_228.INIT = 16'h8000;
LUT4 lut_inst_229 (
  .F(lut_f_229),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_229.INIT = 16'h8000;
LUT4 lut_inst_230 (
  .F(lut_f_230),
  .I0(lut_f_228),
  .I1(lut_f_229),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_230.INIT = 16'h8000;
LUT4 lut_inst_231 (
  .F(lut_f_231),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_231.INIT = 16'h8000;
LUT4 lut_inst_232 (
  .F(lut_f_232),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_232.INIT = 16'h8000;
LUT4 lut_inst_233 (
  .F(lut_f_233),
  .I0(lut_f_231),
  .I1(lut_f_232),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_233.INIT = 16'h8000;
LUT4 lut_inst_234 (
  .F(lut_f_234),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_234.INIT = 16'h8000;
LUT4 lut_inst_235 (
  .F(lut_f_235),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_235.INIT = 16'h8000;
LUT4 lut_inst_236 (
  .F(lut_f_236),
  .I0(lut_f_234),
  .I1(lut_f_235),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_236.INIT = 16'h8000;
LUT4 lut_inst_237 (
  .F(lut_f_237),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_237.INIT = 16'h8000;
LUT4 lut_inst_238 (
  .F(lut_f_238),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_238.INIT = 16'h8000;
LUT4 lut_inst_239 (
  .F(lut_f_239),
  .I0(lut_f_237),
  .I1(lut_f_238),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_239.INIT = 16'h8000;
LUT4 lut_inst_240 (
  .F(lut_f_240),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_240.INIT = 16'h8000;
LUT4 lut_inst_241 (
  .F(lut_f_241),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_241.INIT = 16'h8000;
LUT4 lut_inst_242 (
  .F(lut_f_242),
  .I0(lut_f_240),
  .I1(lut_f_241),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_242.INIT = 16'h8000;
LUT4 lut_inst_243 (
  .F(lut_f_243),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_243.INIT = 16'h8000;
LUT4 lut_inst_244 (
  .F(lut_f_244),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_244.INIT = 16'h8000;
LUT4 lut_inst_245 (
  .F(lut_f_245),
  .I0(lut_f_243),
  .I1(lut_f_244),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_245.INIT = 16'h8000;
LUT4 lut_inst_246 (
  .F(lut_f_246),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_246.INIT = 16'h8000;
LUT4 lut_inst_247 (
  .F(lut_f_247),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_247.INIT = 16'h8000;
LUT4 lut_inst_248 (
  .F(lut_f_248),
  .I0(lut_f_246),
  .I1(lut_f_247),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_248.INIT = 16'h8000;
LUT4 lut_inst_249 (
  .F(lut_f_249),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_249.INIT = 16'h8000;
LUT4 lut_inst_250 (
  .F(lut_f_250),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_250.INIT = 16'h8000;
LUT4 lut_inst_251 (
  .F(lut_f_251),
  .I0(lut_f_249),
  .I1(lut_f_250),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_251.INIT = 16'h8000;
LUT4 lut_inst_252 (
  .F(lut_f_252),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_252.INIT = 16'h8000;
LUT4 lut_inst_253 (
  .F(lut_f_253),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_253.INIT = 16'h8000;
LUT4 lut_inst_254 (
  .F(lut_f_254),
  .I0(lut_f_252),
  .I1(lut_f_253),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_254.INIT = 16'h8000;
LUT4 lut_inst_255 (
  .F(lut_f_255),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_255.INIT = 16'h8000;
LUT4 lut_inst_256 (
  .F(lut_f_256),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_256.INIT = 16'h8000;
LUT4 lut_inst_257 (
  .F(lut_f_257),
  .I0(lut_f_255),
  .I1(lut_f_256),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_257.INIT = 16'h8000;
LUT4 lut_inst_258 (
  .F(lut_f_258),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_258.INIT = 16'h8000;
LUT4 lut_inst_259 (
  .F(lut_f_259),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_259.INIT = 16'h8000;
LUT4 lut_inst_260 (
  .F(lut_f_260),
  .I0(lut_f_258),
  .I1(lut_f_259),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_260.INIT = 16'h8000;
LUT4 lut_inst_261 (
  .F(lut_f_261),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_261.INIT = 16'h8000;
LUT4 lut_inst_262 (
  .F(lut_f_262),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_262.INIT = 16'h8000;
LUT4 lut_inst_263 (
  .F(lut_f_263),
  .I0(lut_f_261),
  .I1(lut_f_262),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_263.INIT = 16'h8000;
LUT4 lut_inst_264 (
  .F(lut_f_264),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_264.INIT = 16'h8000;
LUT4 lut_inst_265 (
  .F(lut_f_265),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_265.INIT = 16'h8000;
LUT4 lut_inst_266 (
  .F(lut_f_266),
  .I0(lut_f_264),
  .I1(lut_f_265),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_266.INIT = 16'h8000;
LUT4 lut_inst_267 (
  .F(lut_f_267),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_267.INIT = 16'h8000;
LUT4 lut_inst_268 (
  .F(lut_f_268),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_268.INIT = 16'h8000;
LUT4 lut_inst_269 (
  .F(lut_f_269),
  .I0(lut_f_267),
  .I1(lut_f_268),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_269.INIT = 16'h8000;
LUT4 lut_inst_270 (
  .F(lut_f_270),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_270.INIT = 16'h8000;
LUT4 lut_inst_271 (
  .F(lut_f_271),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_271.INIT = 16'h8000;
LUT4 lut_inst_272 (
  .F(lut_f_272),
  .I0(lut_f_270),
  .I1(lut_f_271),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_272.INIT = 16'h8000;
LUT4 lut_inst_273 (
  .F(lut_f_273),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_273.INIT = 16'h8000;
LUT4 lut_inst_274 (
  .F(lut_f_274),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_274.INIT = 16'h8000;
LUT4 lut_inst_275 (
  .F(lut_f_275),
  .I0(lut_f_273),
  .I1(lut_f_274),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_275.INIT = 16'h8000;
LUT4 lut_inst_276 (
  .F(lut_f_276),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_276.INIT = 16'h8000;
LUT4 lut_inst_277 (
  .F(lut_f_277),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_277.INIT = 16'h8000;
LUT4 lut_inst_278 (
  .F(lut_f_278),
  .I0(lut_f_276),
  .I1(lut_f_277),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_278.INIT = 16'h8000;
LUT4 lut_inst_279 (
  .F(lut_f_279),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_279.INIT = 16'h8000;
LUT4 lut_inst_280 (
  .F(lut_f_280),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_280.INIT = 16'h8000;
LUT4 lut_inst_281 (
  .F(lut_f_281),
  .I0(lut_f_279),
  .I1(lut_f_280),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_281.INIT = 16'h8000;
LUT4 lut_inst_282 (
  .F(lut_f_282),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_282.INIT = 16'h8000;
LUT4 lut_inst_283 (
  .F(lut_f_283),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_283.INIT = 16'h8000;
LUT4 lut_inst_284 (
  .F(lut_f_284),
  .I0(lut_f_282),
  .I1(lut_f_283),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_284.INIT = 16'h8000;
LUT4 lut_inst_285 (
  .F(lut_f_285),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_285.INIT = 16'h8000;
LUT4 lut_inst_286 (
  .F(lut_f_286),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad9_inv),
  .I3(wad[10])
);
defparam lut_inst_286.INIT = 16'h8000;
LUT4 lut_inst_287 (
  .F(lut_f_287),
  .I0(lut_f_285),
  .I1(lut_f_286),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_287.INIT = 16'h8000;
LUT4 lut_inst_288 (
  .F(lut_f_288),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_288.INIT = 16'h8000;
LUT4 lut_inst_289 (
  .F(lut_f_289),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_289.INIT = 16'h8000;
LUT4 lut_inst_290 (
  .F(lut_f_290),
  .I0(lut_f_288),
  .I1(lut_f_289),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_290.INIT = 16'h8000;
LUT4 lut_inst_291 (
  .F(lut_f_291),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_291.INIT = 16'h8000;
LUT4 lut_inst_292 (
  .F(lut_f_292),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_292.INIT = 16'h8000;
LUT4 lut_inst_293 (
  .F(lut_f_293),
  .I0(lut_f_291),
  .I1(lut_f_292),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_293.INIT = 16'h8000;
LUT4 lut_inst_294 (
  .F(lut_f_294),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_294.INIT = 16'h8000;
LUT4 lut_inst_295 (
  .F(lut_f_295),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_295.INIT = 16'h8000;
LUT4 lut_inst_296 (
  .F(lut_f_296),
  .I0(lut_f_294),
  .I1(lut_f_295),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_296.INIT = 16'h8000;
LUT4 lut_inst_297 (
  .F(lut_f_297),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_297.INIT = 16'h8000;
LUT4 lut_inst_298 (
  .F(lut_f_298),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_298.INIT = 16'h8000;
LUT4 lut_inst_299 (
  .F(lut_f_299),
  .I0(lut_f_297),
  .I1(lut_f_298),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_299.INIT = 16'h8000;
LUT4 lut_inst_300 (
  .F(lut_f_300),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_300.INIT = 16'h8000;
LUT4 lut_inst_301 (
  .F(lut_f_301),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_301.INIT = 16'h8000;
LUT4 lut_inst_302 (
  .F(lut_f_302),
  .I0(lut_f_300),
  .I1(lut_f_301),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_302.INIT = 16'h8000;
LUT4 lut_inst_303 (
  .F(lut_f_303),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_303.INIT = 16'h8000;
LUT4 lut_inst_304 (
  .F(lut_f_304),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_304.INIT = 16'h8000;
LUT4 lut_inst_305 (
  .F(lut_f_305),
  .I0(lut_f_303),
  .I1(lut_f_304),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_305.INIT = 16'h8000;
LUT4 lut_inst_306 (
  .F(lut_f_306),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_306.INIT = 16'h8000;
LUT4 lut_inst_307 (
  .F(lut_f_307),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_307.INIT = 16'h8000;
LUT4 lut_inst_308 (
  .F(lut_f_308),
  .I0(lut_f_306),
  .I1(lut_f_307),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_308.INIT = 16'h8000;
LUT4 lut_inst_309 (
  .F(lut_f_309),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_309.INIT = 16'h8000;
LUT4 lut_inst_310 (
  .F(lut_f_310),
  .I0(wad7_inv),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_310.INIT = 16'h8000;
LUT4 lut_inst_311 (
  .F(lut_f_311),
  .I0(lut_f_309),
  .I1(lut_f_310),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_311.INIT = 16'h8000;
LUT4 lut_inst_312 (
  .F(lut_f_312),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_312.INIT = 16'h8000;
LUT4 lut_inst_313 (
  .F(lut_f_313),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_313.INIT = 16'h8000;
LUT4 lut_inst_314 (
  .F(lut_f_314),
  .I0(lut_f_312),
  .I1(lut_f_313),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_314.INIT = 16'h8000;
LUT4 lut_inst_315 (
  .F(lut_f_315),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_315.INIT = 16'h8000;
LUT4 lut_inst_316 (
  .F(lut_f_316),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_316.INIT = 16'h8000;
LUT4 lut_inst_317 (
  .F(lut_f_317),
  .I0(lut_f_315),
  .I1(lut_f_316),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_317.INIT = 16'h8000;
LUT4 lut_inst_318 (
  .F(lut_f_318),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_318.INIT = 16'h8000;
LUT4 lut_inst_319 (
  .F(lut_f_319),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_319.INIT = 16'h8000;
LUT4 lut_inst_320 (
  .F(lut_f_320),
  .I0(lut_f_318),
  .I1(lut_f_319),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_320.INIT = 16'h8000;
LUT4 lut_inst_321 (
  .F(lut_f_321),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_321.INIT = 16'h8000;
LUT4 lut_inst_322 (
  .F(lut_f_322),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_322.INIT = 16'h8000;
LUT4 lut_inst_323 (
  .F(lut_f_323),
  .I0(lut_f_321),
  .I1(lut_f_322),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_323.INIT = 16'h8000;
LUT4 lut_inst_324 (
  .F(lut_f_324),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_324.INIT = 16'h8000;
LUT4 lut_inst_325 (
  .F(lut_f_325),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_325.INIT = 16'h8000;
LUT4 lut_inst_326 (
  .F(lut_f_326),
  .I0(lut_f_324),
  .I1(lut_f_325),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_326.INIT = 16'h8000;
LUT4 lut_inst_327 (
  .F(lut_f_327),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_327.INIT = 16'h8000;
LUT4 lut_inst_328 (
  .F(lut_f_328),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_328.INIT = 16'h8000;
LUT4 lut_inst_329 (
  .F(lut_f_329),
  .I0(lut_f_327),
  .I1(lut_f_328),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_329.INIT = 16'h8000;
LUT4 lut_inst_330 (
  .F(lut_f_330),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_330.INIT = 16'h8000;
LUT4 lut_inst_331 (
  .F(lut_f_331),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_331.INIT = 16'h8000;
LUT4 lut_inst_332 (
  .F(lut_f_332),
  .I0(lut_f_330),
  .I1(lut_f_331),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_332.INIT = 16'h8000;
LUT4 lut_inst_333 (
  .F(lut_f_333),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_333.INIT = 16'h8000;
LUT4 lut_inst_334 (
  .F(lut_f_334),
  .I0(wad[7]),
  .I1(wad8_inv),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_334.INIT = 16'h8000;
LUT4 lut_inst_335 (
  .F(lut_f_335),
  .I0(lut_f_333),
  .I1(lut_f_334),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_335.INIT = 16'h8000;
LUT4 lut_inst_336 (
  .F(lut_f_336),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_336.INIT = 16'h8000;
LUT4 lut_inst_337 (
  .F(lut_f_337),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_337.INIT = 16'h8000;
LUT4 lut_inst_338 (
  .F(lut_f_338),
  .I0(lut_f_336),
  .I1(lut_f_337),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_338.INIT = 16'h8000;
LUT4 lut_inst_339 (
  .F(lut_f_339),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_339.INIT = 16'h8000;
LUT4 lut_inst_340 (
  .F(lut_f_340),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_340.INIT = 16'h8000;
LUT4 lut_inst_341 (
  .F(lut_f_341),
  .I0(lut_f_339),
  .I1(lut_f_340),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_341.INIT = 16'h8000;
LUT4 lut_inst_342 (
  .F(lut_f_342),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_342.INIT = 16'h8000;
LUT4 lut_inst_343 (
  .F(lut_f_343),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_343.INIT = 16'h8000;
LUT4 lut_inst_344 (
  .F(lut_f_344),
  .I0(lut_f_342),
  .I1(lut_f_343),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_344.INIT = 16'h8000;
LUT4 lut_inst_345 (
  .F(lut_f_345),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_345.INIT = 16'h8000;
LUT4 lut_inst_346 (
  .F(lut_f_346),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_346.INIT = 16'h8000;
LUT4 lut_inst_347 (
  .F(lut_f_347),
  .I0(lut_f_345),
  .I1(lut_f_346),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_347.INIT = 16'h8000;
LUT4 lut_inst_348 (
  .F(lut_f_348),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_348.INIT = 16'h8000;
LUT4 lut_inst_349 (
  .F(lut_f_349),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_349.INIT = 16'h8000;
LUT4 lut_inst_350 (
  .F(lut_f_350),
  .I0(lut_f_348),
  .I1(lut_f_349),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_350.INIT = 16'h8000;
LUT4 lut_inst_351 (
  .F(lut_f_351),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_351.INIT = 16'h8000;
LUT4 lut_inst_352 (
  .F(lut_f_352),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_352.INIT = 16'h8000;
LUT4 lut_inst_353 (
  .F(lut_f_353),
  .I0(lut_f_351),
  .I1(lut_f_352),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_353.INIT = 16'h8000;
LUT4 lut_inst_354 (
  .F(lut_f_354),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_354.INIT = 16'h8000;
LUT4 lut_inst_355 (
  .F(lut_f_355),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_355.INIT = 16'h8000;
LUT4 lut_inst_356 (
  .F(lut_f_356),
  .I0(lut_f_354),
  .I1(lut_f_355),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_356.INIT = 16'h8000;
LUT4 lut_inst_357 (
  .F(lut_f_357),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_357.INIT = 16'h8000;
LUT4 lut_inst_358 (
  .F(lut_f_358),
  .I0(wad7_inv),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_358.INIT = 16'h8000;
LUT4 lut_inst_359 (
  .F(lut_f_359),
  .I0(lut_f_357),
  .I1(lut_f_358),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_359.INIT = 16'h8000;
LUT4 lut_inst_360 (
  .F(lut_f_360),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_360.INIT = 16'h8000;
LUT4 lut_inst_361 (
  .F(lut_f_361),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_361.INIT = 16'h8000;
LUT4 lut_inst_362 (
  .F(lut_f_362),
  .I0(lut_f_360),
  .I1(lut_f_361),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_362.INIT = 16'h8000;
LUT4 lut_inst_363 (
  .F(lut_f_363),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_363.INIT = 16'h8000;
LUT4 lut_inst_364 (
  .F(lut_f_364),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_364.INIT = 16'h8000;
LUT4 lut_inst_365 (
  .F(lut_f_365),
  .I0(lut_f_363),
  .I1(lut_f_364),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_365.INIT = 16'h8000;
LUT4 lut_inst_366 (
  .F(lut_f_366),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_366.INIT = 16'h8000;
LUT4 lut_inst_367 (
  .F(lut_f_367),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_367.INIT = 16'h8000;
LUT4 lut_inst_368 (
  .F(lut_f_368),
  .I0(lut_f_366),
  .I1(lut_f_367),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_368.INIT = 16'h8000;
LUT4 lut_inst_369 (
  .F(lut_f_369),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_369.INIT = 16'h8000;
LUT4 lut_inst_370 (
  .F(lut_f_370),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_370.INIT = 16'h8000;
LUT4 lut_inst_371 (
  .F(lut_f_371),
  .I0(lut_f_369),
  .I1(lut_f_370),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_371.INIT = 16'h8000;
LUT4 lut_inst_372 (
  .F(lut_f_372),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_372.INIT = 16'h8000;
LUT4 lut_inst_373 (
  .F(lut_f_373),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_373.INIT = 16'h8000;
LUT4 lut_inst_374 (
  .F(lut_f_374),
  .I0(lut_f_372),
  .I1(lut_f_373),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_374.INIT = 16'h8000;
LUT4 lut_inst_375 (
  .F(lut_f_375),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_375.INIT = 16'h8000;
LUT4 lut_inst_376 (
  .F(lut_f_376),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_376.INIT = 16'h8000;
LUT4 lut_inst_377 (
  .F(lut_f_377),
  .I0(lut_f_375),
  .I1(lut_f_376),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_377.INIT = 16'h8000;
LUT4 lut_inst_378 (
  .F(lut_f_378),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_378.INIT = 16'h8000;
LUT4 lut_inst_379 (
  .F(lut_f_379),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_379.INIT = 16'h8000;
LUT4 lut_inst_380 (
  .F(lut_f_380),
  .I0(lut_f_378),
  .I1(lut_f_379),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_380.INIT = 16'h8000;
LUT4 lut_inst_381 (
  .F(lut_f_381),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_381.INIT = 16'h8000;
LUT4 lut_inst_382 (
  .F(lut_f_382),
  .I0(wad[7]),
  .I1(wad[8]),
  .I2(wad[9]),
  .I3(wad[10])
);
defparam lut_inst_382.INIT = 16'h8000;
LUT4 lut_inst_383 (
  .F(lut_f_383),
  .I0(lut_f_381),
  .I1(lut_f_382),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_383.INIT = 16'h8000;
RAM16SDP4 ram16sdp_inst_0 (
    .DO(ram16sdp_inst_0_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_2),
    .CLK(clk)
);

defparam ram16sdp_inst_0.INIT_0 = 16'h0000;
defparam ram16sdp_inst_0.INIT_1 = 16'h0000;
defparam ram16sdp_inst_0.INIT_2 = 16'h0000;
defparam ram16sdp_inst_0.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1 (
    .DO(ram16sdp_inst_1_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_2),
    .CLK(clk)
);

defparam ram16sdp_inst_1.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_2 (
    .DO(ram16sdp_inst_2_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_2),
    .CLK(clk)
);

defparam ram16sdp_inst_2.INIT_0 = 16'h0000;
defparam ram16sdp_inst_2.INIT_1 = 16'h0000;
defparam ram16sdp_inst_2.INIT_2 = 16'h0000;
defparam ram16sdp_inst_2.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_3 (
    .DO(ram16sdp_inst_3_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_2),
    .CLK(clk)
);

defparam ram16sdp_inst_3.INIT_0 = 16'h0000;
defparam ram16sdp_inst_3.INIT_1 = 16'h0000;
defparam ram16sdp_inst_3.INIT_2 = 16'h0000;
defparam ram16sdp_inst_3.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_4 (
    .DO(ram16sdp_inst_4_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_2),
    .CLK(clk)
);

defparam ram16sdp_inst_4.INIT_0 = 16'h0000;
defparam ram16sdp_inst_4.INIT_1 = 16'h0000;
defparam ram16sdp_inst_4.INIT_2 = 16'h0000;
defparam ram16sdp_inst_4.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_5 (
    .DO(ram16sdp_inst_5_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_2),
    .CLK(clk)
);

defparam ram16sdp_inst_5.INIT_0 = 16'h0000;
defparam ram16sdp_inst_5.INIT_1 = 16'h0000;
defparam ram16sdp_inst_5.INIT_2 = 16'h0000;
defparam ram16sdp_inst_5.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_6 (
    .DO(ram16sdp_inst_6_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_2),
    .CLK(clk)
);

defparam ram16sdp_inst_6.INIT_0 = 16'h0000;
defparam ram16sdp_inst_6.INIT_1 = 16'h0000;
defparam ram16sdp_inst_6.INIT_2 = 16'h0000;
defparam ram16sdp_inst_6.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_7 (
    .DO(ram16sdp_inst_7_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_2),
    .CLK(clk)
);

defparam ram16sdp_inst_7.INIT_0 = 16'h0000;
defparam ram16sdp_inst_7.INIT_1 = 16'h0000;
defparam ram16sdp_inst_7.INIT_2 = 16'h0000;
defparam ram16sdp_inst_7.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_8 (
    .DO(ram16sdp_inst_8_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_8.INIT_0 = 16'h0000;
defparam ram16sdp_inst_8.INIT_1 = 16'h0000;
defparam ram16sdp_inst_8.INIT_2 = 16'h0000;
defparam ram16sdp_inst_8.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_9 (
    .DO(ram16sdp_inst_9_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_9.INIT_0 = 16'h0000;
defparam ram16sdp_inst_9.INIT_1 = 16'h0000;
defparam ram16sdp_inst_9.INIT_2 = 16'h0000;
defparam ram16sdp_inst_9.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_10 (
    .DO(ram16sdp_inst_10_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_10.INIT_0 = 16'h0000;
defparam ram16sdp_inst_10.INIT_1 = 16'h0000;
defparam ram16sdp_inst_10.INIT_2 = 16'h0000;
defparam ram16sdp_inst_10.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_11 (
    .DO(ram16sdp_inst_11_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_11.INIT_0 = 16'h0000;
defparam ram16sdp_inst_11.INIT_1 = 16'h0000;
defparam ram16sdp_inst_11.INIT_2 = 16'h0000;
defparam ram16sdp_inst_11.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_12 (
    .DO(ram16sdp_inst_12_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_12.INIT_0 = 16'h0000;
defparam ram16sdp_inst_12.INIT_1 = 16'h0000;
defparam ram16sdp_inst_12.INIT_2 = 16'h0000;
defparam ram16sdp_inst_12.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_13 (
    .DO(ram16sdp_inst_13_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_13.INIT_0 = 16'h0000;
defparam ram16sdp_inst_13.INIT_1 = 16'h0000;
defparam ram16sdp_inst_13.INIT_2 = 16'h0000;
defparam ram16sdp_inst_13.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_14 (
    .DO(ram16sdp_inst_14_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_14.INIT_0 = 16'h0000;
defparam ram16sdp_inst_14.INIT_1 = 16'h0000;
defparam ram16sdp_inst_14.INIT_2 = 16'h0000;
defparam ram16sdp_inst_14.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_15 (
    .DO(ram16sdp_inst_15_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_15.INIT_0 = 16'h0000;
defparam ram16sdp_inst_15.INIT_1 = 16'h0000;
defparam ram16sdp_inst_15.INIT_2 = 16'h0000;
defparam ram16sdp_inst_15.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_16 (
    .DO(ram16sdp_inst_16_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_8),
    .CLK(clk)
);

defparam ram16sdp_inst_16.INIT_0 = 16'h0000;
defparam ram16sdp_inst_16.INIT_1 = 16'h0000;
defparam ram16sdp_inst_16.INIT_2 = 16'h0000;
defparam ram16sdp_inst_16.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_17 (
    .DO(ram16sdp_inst_17_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_8),
    .CLK(clk)
);

defparam ram16sdp_inst_17.INIT_0 = 16'h0000;
defparam ram16sdp_inst_17.INIT_1 = 16'h0000;
defparam ram16sdp_inst_17.INIT_2 = 16'h0000;
defparam ram16sdp_inst_17.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_18 (
    .DO(ram16sdp_inst_18_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_8),
    .CLK(clk)
);

defparam ram16sdp_inst_18.INIT_0 = 16'h0000;
defparam ram16sdp_inst_18.INIT_1 = 16'h0000;
defparam ram16sdp_inst_18.INIT_2 = 16'h0000;
defparam ram16sdp_inst_18.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_19 (
    .DO(ram16sdp_inst_19_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_8),
    .CLK(clk)
);

defparam ram16sdp_inst_19.INIT_0 = 16'h0000;
defparam ram16sdp_inst_19.INIT_1 = 16'h0000;
defparam ram16sdp_inst_19.INIT_2 = 16'h0000;
defparam ram16sdp_inst_19.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_20 (
    .DO(ram16sdp_inst_20_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_8),
    .CLK(clk)
);

defparam ram16sdp_inst_20.INIT_0 = 16'h0000;
defparam ram16sdp_inst_20.INIT_1 = 16'h0000;
defparam ram16sdp_inst_20.INIT_2 = 16'h0000;
defparam ram16sdp_inst_20.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_21 (
    .DO(ram16sdp_inst_21_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_8),
    .CLK(clk)
);

defparam ram16sdp_inst_21.INIT_0 = 16'h0000;
defparam ram16sdp_inst_21.INIT_1 = 16'h0000;
defparam ram16sdp_inst_21.INIT_2 = 16'h0000;
defparam ram16sdp_inst_21.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_22 (
    .DO(ram16sdp_inst_22_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_8),
    .CLK(clk)
);

defparam ram16sdp_inst_22.INIT_0 = 16'h0000;
defparam ram16sdp_inst_22.INIT_1 = 16'h0000;
defparam ram16sdp_inst_22.INIT_2 = 16'h0000;
defparam ram16sdp_inst_22.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_23 (
    .DO(ram16sdp_inst_23_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_8),
    .CLK(clk)
);

defparam ram16sdp_inst_23.INIT_0 = 16'h0000;
defparam ram16sdp_inst_23.INIT_1 = 16'h0000;
defparam ram16sdp_inst_23.INIT_2 = 16'h0000;
defparam ram16sdp_inst_23.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_24 (
    .DO(ram16sdp_inst_24_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_24.INIT_0 = 16'h0000;
defparam ram16sdp_inst_24.INIT_1 = 16'h0000;
defparam ram16sdp_inst_24.INIT_2 = 16'h0000;
defparam ram16sdp_inst_24.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_25 (
    .DO(ram16sdp_inst_25_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_25.INIT_0 = 16'h0000;
defparam ram16sdp_inst_25.INIT_1 = 16'h0000;
defparam ram16sdp_inst_25.INIT_2 = 16'h0000;
defparam ram16sdp_inst_25.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_26 (
    .DO(ram16sdp_inst_26_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_26.INIT_0 = 16'h0000;
defparam ram16sdp_inst_26.INIT_1 = 16'h0000;
defparam ram16sdp_inst_26.INIT_2 = 16'h0000;
defparam ram16sdp_inst_26.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_27 (
    .DO(ram16sdp_inst_27_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_27.INIT_0 = 16'h0000;
defparam ram16sdp_inst_27.INIT_1 = 16'h0000;
defparam ram16sdp_inst_27.INIT_2 = 16'h0000;
defparam ram16sdp_inst_27.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_28 (
    .DO(ram16sdp_inst_28_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_28.INIT_0 = 16'h0000;
defparam ram16sdp_inst_28.INIT_1 = 16'h0000;
defparam ram16sdp_inst_28.INIT_2 = 16'h0000;
defparam ram16sdp_inst_28.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_29 (
    .DO(ram16sdp_inst_29_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_29.INIT_0 = 16'h0000;
defparam ram16sdp_inst_29.INIT_1 = 16'h0000;
defparam ram16sdp_inst_29.INIT_2 = 16'h0000;
defparam ram16sdp_inst_29.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_30 (
    .DO(ram16sdp_inst_30_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_30.INIT_0 = 16'h0000;
defparam ram16sdp_inst_30.INIT_1 = 16'h0000;
defparam ram16sdp_inst_30.INIT_2 = 16'h0000;
defparam ram16sdp_inst_30.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_31 (
    .DO(ram16sdp_inst_31_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_31.INIT_0 = 16'h0000;
defparam ram16sdp_inst_31.INIT_1 = 16'h0000;
defparam ram16sdp_inst_31.INIT_2 = 16'h0000;
defparam ram16sdp_inst_31.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_32 (
    .DO(ram16sdp_inst_32_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_14),
    .CLK(clk)
);

defparam ram16sdp_inst_32.INIT_0 = 16'h0000;
defparam ram16sdp_inst_32.INIT_1 = 16'h0000;
defparam ram16sdp_inst_32.INIT_2 = 16'h0000;
defparam ram16sdp_inst_32.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_33 (
    .DO(ram16sdp_inst_33_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_14),
    .CLK(clk)
);

defparam ram16sdp_inst_33.INIT_0 = 16'h0000;
defparam ram16sdp_inst_33.INIT_1 = 16'h0000;
defparam ram16sdp_inst_33.INIT_2 = 16'h0000;
defparam ram16sdp_inst_33.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_34 (
    .DO(ram16sdp_inst_34_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_14),
    .CLK(clk)
);

defparam ram16sdp_inst_34.INIT_0 = 16'h0000;
defparam ram16sdp_inst_34.INIT_1 = 16'h0000;
defparam ram16sdp_inst_34.INIT_2 = 16'h0000;
defparam ram16sdp_inst_34.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_35 (
    .DO(ram16sdp_inst_35_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_14),
    .CLK(clk)
);

defparam ram16sdp_inst_35.INIT_0 = 16'h0000;
defparam ram16sdp_inst_35.INIT_1 = 16'h0000;
defparam ram16sdp_inst_35.INIT_2 = 16'h0000;
defparam ram16sdp_inst_35.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_36 (
    .DO(ram16sdp_inst_36_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_14),
    .CLK(clk)
);

defparam ram16sdp_inst_36.INIT_0 = 16'h0000;
defparam ram16sdp_inst_36.INIT_1 = 16'h0000;
defparam ram16sdp_inst_36.INIT_2 = 16'h0000;
defparam ram16sdp_inst_36.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_37 (
    .DO(ram16sdp_inst_37_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_14),
    .CLK(clk)
);

defparam ram16sdp_inst_37.INIT_0 = 16'h0000;
defparam ram16sdp_inst_37.INIT_1 = 16'h0000;
defparam ram16sdp_inst_37.INIT_2 = 16'h0000;
defparam ram16sdp_inst_37.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_38 (
    .DO(ram16sdp_inst_38_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_14),
    .CLK(clk)
);

defparam ram16sdp_inst_38.INIT_0 = 16'h0000;
defparam ram16sdp_inst_38.INIT_1 = 16'h0000;
defparam ram16sdp_inst_38.INIT_2 = 16'h0000;
defparam ram16sdp_inst_38.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_39 (
    .DO(ram16sdp_inst_39_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_14),
    .CLK(clk)
);

defparam ram16sdp_inst_39.INIT_0 = 16'h0000;
defparam ram16sdp_inst_39.INIT_1 = 16'h0000;
defparam ram16sdp_inst_39.INIT_2 = 16'h0000;
defparam ram16sdp_inst_39.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_40 (
    .DO(ram16sdp_inst_40_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_40.INIT_0 = 16'h0000;
defparam ram16sdp_inst_40.INIT_1 = 16'h0000;
defparam ram16sdp_inst_40.INIT_2 = 16'h0000;
defparam ram16sdp_inst_40.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_41 (
    .DO(ram16sdp_inst_41_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_41.INIT_0 = 16'h0000;
defparam ram16sdp_inst_41.INIT_1 = 16'h0000;
defparam ram16sdp_inst_41.INIT_2 = 16'h0000;
defparam ram16sdp_inst_41.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_42 (
    .DO(ram16sdp_inst_42_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_42.INIT_0 = 16'h0000;
defparam ram16sdp_inst_42.INIT_1 = 16'h0000;
defparam ram16sdp_inst_42.INIT_2 = 16'h0000;
defparam ram16sdp_inst_42.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_43 (
    .DO(ram16sdp_inst_43_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_43.INIT_0 = 16'h0000;
defparam ram16sdp_inst_43.INIT_1 = 16'h0000;
defparam ram16sdp_inst_43.INIT_2 = 16'h0000;
defparam ram16sdp_inst_43.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_44 (
    .DO(ram16sdp_inst_44_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_44.INIT_0 = 16'h0000;
defparam ram16sdp_inst_44.INIT_1 = 16'h0000;
defparam ram16sdp_inst_44.INIT_2 = 16'h0000;
defparam ram16sdp_inst_44.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_45 (
    .DO(ram16sdp_inst_45_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_45.INIT_0 = 16'h0000;
defparam ram16sdp_inst_45.INIT_1 = 16'h0000;
defparam ram16sdp_inst_45.INIT_2 = 16'h0000;
defparam ram16sdp_inst_45.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_46 (
    .DO(ram16sdp_inst_46_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_46.INIT_0 = 16'h0000;
defparam ram16sdp_inst_46.INIT_1 = 16'h0000;
defparam ram16sdp_inst_46.INIT_2 = 16'h0000;
defparam ram16sdp_inst_46.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_47 (
    .DO(ram16sdp_inst_47_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_47.INIT_0 = 16'h0000;
defparam ram16sdp_inst_47.INIT_1 = 16'h0000;
defparam ram16sdp_inst_47.INIT_2 = 16'h0000;
defparam ram16sdp_inst_47.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_48 (
    .DO(ram16sdp_inst_48_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_20),
    .CLK(clk)
);

defparam ram16sdp_inst_48.INIT_0 = 16'h0000;
defparam ram16sdp_inst_48.INIT_1 = 16'h0000;
defparam ram16sdp_inst_48.INIT_2 = 16'h0000;
defparam ram16sdp_inst_48.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_49 (
    .DO(ram16sdp_inst_49_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_20),
    .CLK(clk)
);

defparam ram16sdp_inst_49.INIT_0 = 16'h0000;
defparam ram16sdp_inst_49.INIT_1 = 16'h0000;
defparam ram16sdp_inst_49.INIT_2 = 16'h0000;
defparam ram16sdp_inst_49.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_50 (
    .DO(ram16sdp_inst_50_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_20),
    .CLK(clk)
);

defparam ram16sdp_inst_50.INIT_0 = 16'h0000;
defparam ram16sdp_inst_50.INIT_1 = 16'h0000;
defparam ram16sdp_inst_50.INIT_2 = 16'h0000;
defparam ram16sdp_inst_50.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_51 (
    .DO(ram16sdp_inst_51_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_20),
    .CLK(clk)
);

defparam ram16sdp_inst_51.INIT_0 = 16'h0000;
defparam ram16sdp_inst_51.INIT_1 = 16'h0000;
defparam ram16sdp_inst_51.INIT_2 = 16'h0000;
defparam ram16sdp_inst_51.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_52 (
    .DO(ram16sdp_inst_52_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_20),
    .CLK(clk)
);

defparam ram16sdp_inst_52.INIT_0 = 16'h0000;
defparam ram16sdp_inst_52.INIT_1 = 16'h0000;
defparam ram16sdp_inst_52.INIT_2 = 16'h0000;
defparam ram16sdp_inst_52.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_53 (
    .DO(ram16sdp_inst_53_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_20),
    .CLK(clk)
);

defparam ram16sdp_inst_53.INIT_0 = 16'h0000;
defparam ram16sdp_inst_53.INIT_1 = 16'h0000;
defparam ram16sdp_inst_53.INIT_2 = 16'h0000;
defparam ram16sdp_inst_53.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_54 (
    .DO(ram16sdp_inst_54_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_20),
    .CLK(clk)
);

defparam ram16sdp_inst_54.INIT_0 = 16'h0000;
defparam ram16sdp_inst_54.INIT_1 = 16'h0000;
defparam ram16sdp_inst_54.INIT_2 = 16'h0000;
defparam ram16sdp_inst_54.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_55 (
    .DO(ram16sdp_inst_55_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_20),
    .CLK(clk)
);

defparam ram16sdp_inst_55.INIT_0 = 16'h0000;
defparam ram16sdp_inst_55.INIT_1 = 16'h0000;
defparam ram16sdp_inst_55.INIT_2 = 16'h0000;
defparam ram16sdp_inst_55.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_56 (
    .DO(ram16sdp_inst_56_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_56.INIT_0 = 16'h0000;
defparam ram16sdp_inst_56.INIT_1 = 16'h0000;
defparam ram16sdp_inst_56.INIT_2 = 16'h0000;
defparam ram16sdp_inst_56.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_57 (
    .DO(ram16sdp_inst_57_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_57.INIT_0 = 16'h0000;
defparam ram16sdp_inst_57.INIT_1 = 16'h0000;
defparam ram16sdp_inst_57.INIT_2 = 16'h0000;
defparam ram16sdp_inst_57.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_58 (
    .DO(ram16sdp_inst_58_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_58.INIT_0 = 16'h0000;
defparam ram16sdp_inst_58.INIT_1 = 16'h0000;
defparam ram16sdp_inst_58.INIT_2 = 16'h0000;
defparam ram16sdp_inst_58.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_59 (
    .DO(ram16sdp_inst_59_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_59.INIT_0 = 16'h0000;
defparam ram16sdp_inst_59.INIT_1 = 16'h0000;
defparam ram16sdp_inst_59.INIT_2 = 16'h0000;
defparam ram16sdp_inst_59.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_60 (
    .DO(ram16sdp_inst_60_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_60.INIT_0 = 16'h0000;
defparam ram16sdp_inst_60.INIT_1 = 16'h0000;
defparam ram16sdp_inst_60.INIT_2 = 16'h0000;
defparam ram16sdp_inst_60.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_61 (
    .DO(ram16sdp_inst_61_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_61.INIT_0 = 16'h0000;
defparam ram16sdp_inst_61.INIT_1 = 16'h0000;
defparam ram16sdp_inst_61.INIT_2 = 16'h0000;
defparam ram16sdp_inst_61.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_62 (
    .DO(ram16sdp_inst_62_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_62.INIT_0 = 16'h0000;
defparam ram16sdp_inst_62.INIT_1 = 16'h0000;
defparam ram16sdp_inst_62.INIT_2 = 16'h0000;
defparam ram16sdp_inst_62.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_63 (
    .DO(ram16sdp_inst_63_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_63.INIT_0 = 16'h0000;
defparam ram16sdp_inst_63.INIT_1 = 16'h0000;
defparam ram16sdp_inst_63.INIT_2 = 16'h0000;
defparam ram16sdp_inst_63.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_64 (
    .DO(ram16sdp_inst_64_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_26),
    .CLK(clk)
);

defparam ram16sdp_inst_64.INIT_0 = 16'h0000;
defparam ram16sdp_inst_64.INIT_1 = 16'h0000;
defparam ram16sdp_inst_64.INIT_2 = 16'h0000;
defparam ram16sdp_inst_64.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_65 (
    .DO(ram16sdp_inst_65_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_26),
    .CLK(clk)
);

defparam ram16sdp_inst_65.INIT_0 = 16'h0000;
defparam ram16sdp_inst_65.INIT_1 = 16'h0000;
defparam ram16sdp_inst_65.INIT_2 = 16'h0000;
defparam ram16sdp_inst_65.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_66 (
    .DO(ram16sdp_inst_66_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_26),
    .CLK(clk)
);

defparam ram16sdp_inst_66.INIT_0 = 16'h0000;
defparam ram16sdp_inst_66.INIT_1 = 16'h0000;
defparam ram16sdp_inst_66.INIT_2 = 16'h0000;
defparam ram16sdp_inst_66.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_67 (
    .DO(ram16sdp_inst_67_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_26),
    .CLK(clk)
);

defparam ram16sdp_inst_67.INIT_0 = 16'h0000;
defparam ram16sdp_inst_67.INIT_1 = 16'h0000;
defparam ram16sdp_inst_67.INIT_2 = 16'h0000;
defparam ram16sdp_inst_67.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_68 (
    .DO(ram16sdp_inst_68_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_26),
    .CLK(clk)
);

defparam ram16sdp_inst_68.INIT_0 = 16'h0000;
defparam ram16sdp_inst_68.INIT_1 = 16'h0000;
defparam ram16sdp_inst_68.INIT_2 = 16'h0000;
defparam ram16sdp_inst_68.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_69 (
    .DO(ram16sdp_inst_69_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_26),
    .CLK(clk)
);

defparam ram16sdp_inst_69.INIT_0 = 16'h0000;
defparam ram16sdp_inst_69.INIT_1 = 16'h0000;
defparam ram16sdp_inst_69.INIT_2 = 16'h0000;
defparam ram16sdp_inst_69.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_70 (
    .DO(ram16sdp_inst_70_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_26),
    .CLK(clk)
);

defparam ram16sdp_inst_70.INIT_0 = 16'h0000;
defparam ram16sdp_inst_70.INIT_1 = 16'h0000;
defparam ram16sdp_inst_70.INIT_2 = 16'h0000;
defparam ram16sdp_inst_70.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_71 (
    .DO(ram16sdp_inst_71_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_26),
    .CLK(clk)
);

defparam ram16sdp_inst_71.INIT_0 = 16'h0000;
defparam ram16sdp_inst_71.INIT_1 = 16'h0000;
defparam ram16sdp_inst_71.INIT_2 = 16'h0000;
defparam ram16sdp_inst_71.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_72 (
    .DO(ram16sdp_inst_72_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_72.INIT_0 = 16'h0000;
defparam ram16sdp_inst_72.INIT_1 = 16'h0000;
defparam ram16sdp_inst_72.INIT_2 = 16'h0000;
defparam ram16sdp_inst_72.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_73 (
    .DO(ram16sdp_inst_73_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_73.INIT_0 = 16'h0000;
defparam ram16sdp_inst_73.INIT_1 = 16'h0000;
defparam ram16sdp_inst_73.INIT_2 = 16'h0000;
defparam ram16sdp_inst_73.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_74 (
    .DO(ram16sdp_inst_74_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_74.INIT_0 = 16'h0000;
defparam ram16sdp_inst_74.INIT_1 = 16'h0000;
defparam ram16sdp_inst_74.INIT_2 = 16'h0000;
defparam ram16sdp_inst_74.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_75 (
    .DO(ram16sdp_inst_75_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_75.INIT_0 = 16'h0000;
defparam ram16sdp_inst_75.INIT_1 = 16'h0000;
defparam ram16sdp_inst_75.INIT_2 = 16'h0000;
defparam ram16sdp_inst_75.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_76 (
    .DO(ram16sdp_inst_76_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_76.INIT_0 = 16'h0000;
defparam ram16sdp_inst_76.INIT_1 = 16'h0000;
defparam ram16sdp_inst_76.INIT_2 = 16'h0000;
defparam ram16sdp_inst_76.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_77 (
    .DO(ram16sdp_inst_77_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_77.INIT_0 = 16'h0000;
defparam ram16sdp_inst_77.INIT_1 = 16'h0000;
defparam ram16sdp_inst_77.INIT_2 = 16'h0000;
defparam ram16sdp_inst_77.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_78 (
    .DO(ram16sdp_inst_78_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_78.INIT_0 = 16'h0000;
defparam ram16sdp_inst_78.INIT_1 = 16'h0000;
defparam ram16sdp_inst_78.INIT_2 = 16'h0000;
defparam ram16sdp_inst_78.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_79 (
    .DO(ram16sdp_inst_79_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_79.INIT_0 = 16'h0000;
defparam ram16sdp_inst_79.INIT_1 = 16'h0000;
defparam ram16sdp_inst_79.INIT_2 = 16'h0000;
defparam ram16sdp_inst_79.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_80 (
    .DO(ram16sdp_inst_80_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_32),
    .CLK(clk)
);

defparam ram16sdp_inst_80.INIT_0 = 16'h0000;
defparam ram16sdp_inst_80.INIT_1 = 16'h0000;
defparam ram16sdp_inst_80.INIT_2 = 16'h0000;
defparam ram16sdp_inst_80.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_81 (
    .DO(ram16sdp_inst_81_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_32),
    .CLK(clk)
);

defparam ram16sdp_inst_81.INIT_0 = 16'h0000;
defparam ram16sdp_inst_81.INIT_1 = 16'h0000;
defparam ram16sdp_inst_81.INIT_2 = 16'h0000;
defparam ram16sdp_inst_81.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_82 (
    .DO(ram16sdp_inst_82_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_32),
    .CLK(clk)
);

defparam ram16sdp_inst_82.INIT_0 = 16'h0000;
defparam ram16sdp_inst_82.INIT_1 = 16'h0000;
defparam ram16sdp_inst_82.INIT_2 = 16'h0000;
defparam ram16sdp_inst_82.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_83 (
    .DO(ram16sdp_inst_83_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_32),
    .CLK(clk)
);

defparam ram16sdp_inst_83.INIT_0 = 16'h0000;
defparam ram16sdp_inst_83.INIT_1 = 16'h0000;
defparam ram16sdp_inst_83.INIT_2 = 16'h0000;
defparam ram16sdp_inst_83.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_84 (
    .DO(ram16sdp_inst_84_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_32),
    .CLK(clk)
);

defparam ram16sdp_inst_84.INIT_0 = 16'h0000;
defparam ram16sdp_inst_84.INIT_1 = 16'h0000;
defparam ram16sdp_inst_84.INIT_2 = 16'h0000;
defparam ram16sdp_inst_84.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_85 (
    .DO(ram16sdp_inst_85_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_32),
    .CLK(clk)
);

defparam ram16sdp_inst_85.INIT_0 = 16'h0000;
defparam ram16sdp_inst_85.INIT_1 = 16'h0000;
defparam ram16sdp_inst_85.INIT_2 = 16'h0000;
defparam ram16sdp_inst_85.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_86 (
    .DO(ram16sdp_inst_86_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_32),
    .CLK(clk)
);

defparam ram16sdp_inst_86.INIT_0 = 16'h0000;
defparam ram16sdp_inst_86.INIT_1 = 16'h0000;
defparam ram16sdp_inst_86.INIT_2 = 16'h0000;
defparam ram16sdp_inst_86.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_87 (
    .DO(ram16sdp_inst_87_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_32),
    .CLK(clk)
);

defparam ram16sdp_inst_87.INIT_0 = 16'h0000;
defparam ram16sdp_inst_87.INIT_1 = 16'h0000;
defparam ram16sdp_inst_87.INIT_2 = 16'h0000;
defparam ram16sdp_inst_87.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_88 (
    .DO(ram16sdp_inst_88_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_88.INIT_0 = 16'h0000;
defparam ram16sdp_inst_88.INIT_1 = 16'h0000;
defparam ram16sdp_inst_88.INIT_2 = 16'h0000;
defparam ram16sdp_inst_88.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_89 (
    .DO(ram16sdp_inst_89_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_89.INIT_0 = 16'h0000;
defparam ram16sdp_inst_89.INIT_1 = 16'h0000;
defparam ram16sdp_inst_89.INIT_2 = 16'h0000;
defparam ram16sdp_inst_89.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_90 (
    .DO(ram16sdp_inst_90_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_90.INIT_0 = 16'h0000;
defparam ram16sdp_inst_90.INIT_1 = 16'h0000;
defparam ram16sdp_inst_90.INIT_2 = 16'h0000;
defparam ram16sdp_inst_90.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_91 (
    .DO(ram16sdp_inst_91_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_91.INIT_0 = 16'h0000;
defparam ram16sdp_inst_91.INIT_1 = 16'h0000;
defparam ram16sdp_inst_91.INIT_2 = 16'h0000;
defparam ram16sdp_inst_91.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_92 (
    .DO(ram16sdp_inst_92_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_92.INIT_0 = 16'h0000;
defparam ram16sdp_inst_92.INIT_1 = 16'h0000;
defparam ram16sdp_inst_92.INIT_2 = 16'h0000;
defparam ram16sdp_inst_92.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_93 (
    .DO(ram16sdp_inst_93_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_93.INIT_0 = 16'h0000;
defparam ram16sdp_inst_93.INIT_1 = 16'h0000;
defparam ram16sdp_inst_93.INIT_2 = 16'h0000;
defparam ram16sdp_inst_93.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_94 (
    .DO(ram16sdp_inst_94_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_94.INIT_0 = 16'h0000;
defparam ram16sdp_inst_94.INIT_1 = 16'h0000;
defparam ram16sdp_inst_94.INIT_2 = 16'h0000;
defparam ram16sdp_inst_94.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_95 (
    .DO(ram16sdp_inst_95_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_95.INIT_0 = 16'h0000;
defparam ram16sdp_inst_95.INIT_1 = 16'h0000;
defparam ram16sdp_inst_95.INIT_2 = 16'h0000;
defparam ram16sdp_inst_95.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_96 (
    .DO(ram16sdp_inst_96_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_38),
    .CLK(clk)
);

defparam ram16sdp_inst_96.INIT_0 = 16'h0000;
defparam ram16sdp_inst_96.INIT_1 = 16'h0000;
defparam ram16sdp_inst_96.INIT_2 = 16'h0000;
defparam ram16sdp_inst_96.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_97 (
    .DO(ram16sdp_inst_97_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_38),
    .CLK(clk)
);

defparam ram16sdp_inst_97.INIT_0 = 16'h0000;
defparam ram16sdp_inst_97.INIT_1 = 16'h0000;
defparam ram16sdp_inst_97.INIT_2 = 16'h0000;
defparam ram16sdp_inst_97.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_98 (
    .DO(ram16sdp_inst_98_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_38),
    .CLK(clk)
);

defparam ram16sdp_inst_98.INIT_0 = 16'h0000;
defparam ram16sdp_inst_98.INIT_1 = 16'h0000;
defparam ram16sdp_inst_98.INIT_2 = 16'h0000;
defparam ram16sdp_inst_98.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_99 (
    .DO(ram16sdp_inst_99_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_38),
    .CLK(clk)
);

defparam ram16sdp_inst_99.INIT_0 = 16'h0000;
defparam ram16sdp_inst_99.INIT_1 = 16'h0000;
defparam ram16sdp_inst_99.INIT_2 = 16'h0000;
defparam ram16sdp_inst_99.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_100 (
    .DO(ram16sdp_inst_100_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_38),
    .CLK(clk)
);

defparam ram16sdp_inst_100.INIT_0 = 16'h0000;
defparam ram16sdp_inst_100.INIT_1 = 16'h0000;
defparam ram16sdp_inst_100.INIT_2 = 16'h0000;
defparam ram16sdp_inst_100.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_101 (
    .DO(ram16sdp_inst_101_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_38),
    .CLK(clk)
);

defparam ram16sdp_inst_101.INIT_0 = 16'h0000;
defparam ram16sdp_inst_101.INIT_1 = 16'h0000;
defparam ram16sdp_inst_101.INIT_2 = 16'h0000;
defparam ram16sdp_inst_101.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_102 (
    .DO(ram16sdp_inst_102_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_38),
    .CLK(clk)
);

defparam ram16sdp_inst_102.INIT_0 = 16'h0000;
defparam ram16sdp_inst_102.INIT_1 = 16'h0000;
defparam ram16sdp_inst_102.INIT_2 = 16'h0000;
defparam ram16sdp_inst_102.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_103 (
    .DO(ram16sdp_inst_103_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_38),
    .CLK(clk)
);

defparam ram16sdp_inst_103.INIT_0 = 16'h0000;
defparam ram16sdp_inst_103.INIT_1 = 16'h0000;
defparam ram16sdp_inst_103.INIT_2 = 16'h0000;
defparam ram16sdp_inst_103.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_104 (
    .DO(ram16sdp_inst_104_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_104.INIT_0 = 16'h0000;
defparam ram16sdp_inst_104.INIT_1 = 16'h0000;
defparam ram16sdp_inst_104.INIT_2 = 16'h0000;
defparam ram16sdp_inst_104.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_105 (
    .DO(ram16sdp_inst_105_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_105.INIT_0 = 16'h0000;
defparam ram16sdp_inst_105.INIT_1 = 16'h0000;
defparam ram16sdp_inst_105.INIT_2 = 16'h0000;
defparam ram16sdp_inst_105.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_106 (
    .DO(ram16sdp_inst_106_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_106.INIT_0 = 16'h0000;
defparam ram16sdp_inst_106.INIT_1 = 16'h0000;
defparam ram16sdp_inst_106.INIT_2 = 16'h0000;
defparam ram16sdp_inst_106.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_107 (
    .DO(ram16sdp_inst_107_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_107.INIT_0 = 16'h0000;
defparam ram16sdp_inst_107.INIT_1 = 16'h0000;
defparam ram16sdp_inst_107.INIT_2 = 16'h0000;
defparam ram16sdp_inst_107.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_108 (
    .DO(ram16sdp_inst_108_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_108.INIT_0 = 16'h0000;
defparam ram16sdp_inst_108.INIT_1 = 16'h0000;
defparam ram16sdp_inst_108.INIT_2 = 16'h0000;
defparam ram16sdp_inst_108.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_109 (
    .DO(ram16sdp_inst_109_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_109.INIT_0 = 16'h0000;
defparam ram16sdp_inst_109.INIT_1 = 16'h0000;
defparam ram16sdp_inst_109.INIT_2 = 16'h0000;
defparam ram16sdp_inst_109.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_110 (
    .DO(ram16sdp_inst_110_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_110.INIT_0 = 16'h0000;
defparam ram16sdp_inst_110.INIT_1 = 16'h0000;
defparam ram16sdp_inst_110.INIT_2 = 16'h0000;
defparam ram16sdp_inst_110.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_111 (
    .DO(ram16sdp_inst_111_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_111.INIT_0 = 16'h0000;
defparam ram16sdp_inst_111.INIT_1 = 16'h0000;
defparam ram16sdp_inst_111.INIT_2 = 16'h0000;
defparam ram16sdp_inst_111.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_112 (
    .DO(ram16sdp_inst_112_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_44),
    .CLK(clk)
);

defparam ram16sdp_inst_112.INIT_0 = 16'h0000;
defparam ram16sdp_inst_112.INIT_1 = 16'h0000;
defparam ram16sdp_inst_112.INIT_2 = 16'h0000;
defparam ram16sdp_inst_112.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_113 (
    .DO(ram16sdp_inst_113_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_44),
    .CLK(clk)
);

defparam ram16sdp_inst_113.INIT_0 = 16'h0000;
defparam ram16sdp_inst_113.INIT_1 = 16'h0000;
defparam ram16sdp_inst_113.INIT_2 = 16'h0000;
defparam ram16sdp_inst_113.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_114 (
    .DO(ram16sdp_inst_114_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_44),
    .CLK(clk)
);

defparam ram16sdp_inst_114.INIT_0 = 16'h0000;
defparam ram16sdp_inst_114.INIT_1 = 16'h0000;
defparam ram16sdp_inst_114.INIT_2 = 16'h0000;
defparam ram16sdp_inst_114.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_115 (
    .DO(ram16sdp_inst_115_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_44),
    .CLK(clk)
);

defparam ram16sdp_inst_115.INIT_0 = 16'h0000;
defparam ram16sdp_inst_115.INIT_1 = 16'h0000;
defparam ram16sdp_inst_115.INIT_2 = 16'h0000;
defparam ram16sdp_inst_115.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_116 (
    .DO(ram16sdp_inst_116_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_44),
    .CLK(clk)
);

defparam ram16sdp_inst_116.INIT_0 = 16'h0000;
defparam ram16sdp_inst_116.INIT_1 = 16'h0000;
defparam ram16sdp_inst_116.INIT_2 = 16'h0000;
defparam ram16sdp_inst_116.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_117 (
    .DO(ram16sdp_inst_117_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_44),
    .CLK(clk)
);

defparam ram16sdp_inst_117.INIT_0 = 16'h0000;
defparam ram16sdp_inst_117.INIT_1 = 16'h0000;
defparam ram16sdp_inst_117.INIT_2 = 16'h0000;
defparam ram16sdp_inst_117.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_118 (
    .DO(ram16sdp_inst_118_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_44),
    .CLK(clk)
);

defparam ram16sdp_inst_118.INIT_0 = 16'h0000;
defparam ram16sdp_inst_118.INIT_1 = 16'h0000;
defparam ram16sdp_inst_118.INIT_2 = 16'h0000;
defparam ram16sdp_inst_118.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_119 (
    .DO(ram16sdp_inst_119_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_44),
    .CLK(clk)
);

defparam ram16sdp_inst_119.INIT_0 = 16'h0000;
defparam ram16sdp_inst_119.INIT_1 = 16'h0000;
defparam ram16sdp_inst_119.INIT_2 = 16'h0000;
defparam ram16sdp_inst_119.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_120 (
    .DO(ram16sdp_inst_120_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_120.INIT_0 = 16'h0000;
defparam ram16sdp_inst_120.INIT_1 = 16'h0000;
defparam ram16sdp_inst_120.INIT_2 = 16'h0000;
defparam ram16sdp_inst_120.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_121 (
    .DO(ram16sdp_inst_121_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_121.INIT_0 = 16'h0000;
defparam ram16sdp_inst_121.INIT_1 = 16'h0000;
defparam ram16sdp_inst_121.INIT_2 = 16'h0000;
defparam ram16sdp_inst_121.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_122 (
    .DO(ram16sdp_inst_122_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_122.INIT_0 = 16'h0000;
defparam ram16sdp_inst_122.INIT_1 = 16'h0000;
defparam ram16sdp_inst_122.INIT_2 = 16'h0000;
defparam ram16sdp_inst_122.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_123 (
    .DO(ram16sdp_inst_123_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_123.INIT_0 = 16'h0000;
defparam ram16sdp_inst_123.INIT_1 = 16'h0000;
defparam ram16sdp_inst_123.INIT_2 = 16'h0000;
defparam ram16sdp_inst_123.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_124 (
    .DO(ram16sdp_inst_124_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_124.INIT_0 = 16'h0000;
defparam ram16sdp_inst_124.INIT_1 = 16'h0000;
defparam ram16sdp_inst_124.INIT_2 = 16'h0000;
defparam ram16sdp_inst_124.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_125 (
    .DO(ram16sdp_inst_125_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_125.INIT_0 = 16'h0000;
defparam ram16sdp_inst_125.INIT_1 = 16'h0000;
defparam ram16sdp_inst_125.INIT_2 = 16'h0000;
defparam ram16sdp_inst_125.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_126 (
    .DO(ram16sdp_inst_126_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_126.INIT_0 = 16'h0000;
defparam ram16sdp_inst_126.INIT_1 = 16'h0000;
defparam ram16sdp_inst_126.INIT_2 = 16'h0000;
defparam ram16sdp_inst_126.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_127 (
    .DO(ram16sdp_inst_127_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_127.INIT_0 = 16'h0000;
defparam ram16sdp_inst_127.INIT_1 = 16'h0000;
defparam ram16sdp_inst_127.INIT_2 = 16'h0000;
defparam ram16sdp_inst_127.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_128 (
    .DO(ram16sdp_inst_128_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_50),
    .CLK(clk)
);

defparam ram16sdp_inst_128.INIT_0 = 16'h0000;
defparam ram16sdp_inst_128.INIT_1 = 16'h0000;
defparam ram16sdp_inst_128.INIT_2 = 16'h0000;
defparam ram16sdp_inst_128.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_129 (
    .DO(ram16sdp_inst_129_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_50),
    .CLK(clk)
);

defparam ram16sdp_inst_129.INIT_0 = 16'h0000;
defparam ram16sdp_inst_129.INIT_1 = 16'h0000;
defparam ram16sdp_inst_129.INIT_2 = 16'h0000;
defparam ram16sdp_inst_129.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_130 (
    .DO(ram16sdp_inst_130_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_50),
    .CLK(clk)
);

defparam ram16sdp_inst_130.INIT_0 = 16'h0000;
defparam ram16sdp_inst_130.INIT_1 = 16'h0000;
defparam ram16sdp_inst_130.INIT_2 = 16'h0000;
defparam ram16sdp_inst_130.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_131 (
    .DO(ram16sdp_inst_131_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_50),
    .CLK(clk)
);

defparam ram16sdp_inst_131.INIT_0 = 16'h0000;
defparam ram16sdp_inst_131.INIT_1 = 16'h0000;
defparam ram16sdp_inst_131.INIT_2 = 16'h0000;
defparam ram16sdp_inst_131.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_132 (
    .DO(ram16sdp_inst_132_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_50),
    .CLK(clk)
);

defparam ram16sdp_inst_132.INIT_0 = 16'h0000;
defparam ram16sdp_inst_132.INIT_1 = 16'h0000;
defparam ram16sdp_inst_132.INIT_2 = 16'h0000;
defparam ram16sdp_inst_132.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_133 (
    .DO(ram16sdp_inst_133_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_50),
    .CLK(clk)
);

defparam ram16sdp_inst_133.INIT_0 = 16'h0000;
defparam ram16sdp_inst_133.INIT_1 = 16'h0000;
defparam ram16sdp_inst_133.INIT_2 = 16'h0000;
defparam ram16sdp_inst_133.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_134 (
    .DO(ram16sdp_inst_134_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_50),
    .CLK(clk)
);

defparam ram16sdp_inst_134.INIT_0 = 16'h0000;
defparam ram16sdp_inst_134.INIT_1 = 16'h0000;
defparam ram16sdp_inst_134.INIT_2 = 16'h0000;
defparam ram16sdp_inst_134.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_135 (
    .DO(ram16sdp_inst_135_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_50),
    .CLK(clk)
);

defparam ram16sdp_inst_135.INIT_0 = 16'h0000;
defparam ram16sdp_inst_135.INIT_1 = 16'h0000;
defparam ram16sdp_inst_135.INIT_2 = 16'h0000;
defparam ram16sdp_inst_135.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_136 (
    .DO(ram16sdp_inst_136_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_136.INIT_0 = 16'h0000;
defparam ram16sdp_inst_136.INIT_1 = 16'h0000;
defparam ram16sdp_inst_136.INIT_2 = 16'h0000;
defparam ram16sdp_inst_136.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_137 (
    .DO(ram16sdp_inst_137_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_137.INIT_0 = 16'h0000;
defparam ram16sdp_inst_137.INIT_1 = 16'h0000;
defparam ram16sdp_inst_137.INIT_2 = 16'h0000;
defparam ram16sdp_inst_137.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_138 (
    .DO(ram16sdp_inst_138_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_138.INIT_0 = 16'h0000;
defparam ram16sdp_inst_138.INIT_1 = 16'h0000;
defparam ram16sdp_inst_138.INIT_2 = 16'h0000;
defparam ram16sdp_inst_138.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_139 (
    .DO(ram16sdp_inst_139_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_139.INIT_0 = 16'h0000;
defparam ram16sdp_inst_139.INIT_1 = 16'h0000;
defparam ram16sdp_inst_139.INIT_2 = 16'h0000;
defparam ram16sdp_inst_139.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_140 (
    .DO(ram16sdp_inst_140_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_140.INIT_0 = 16'h0000;
defparam ram16sdp_inst_140.INIT_1 = 16'h0000;
defparam ram16sdp_inst_140.INIT_2 = 16'h0000;
defparam ram16sdp_inst_140.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_141 (
    .DO(ram16sdp_inst_141_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_141.INIT_0 = 16'h0000;
defparam ram16sdp_inst_141.INIT_1 = 16'h0000;
defparam ram16sdp_inst_141.INIT_2 = 16'h0000;
defparam ram16sdp_inst_141.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_142 (
    .DO(ram16sdp_inst_142_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_142.INIT_0 = 16'h0000;
defparam ram16sdp_inst_142.INIT_1 = 16'h0000;
defparam ram16sdp_inst_142.INIT_2 = 16'h0000;
defparam ram16sdp_inst_142.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_143 (
    .DO(ram16sdp_inst_143_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_143.INIT_0 = 16'h0000;
defparam ram16sdp_inst_143.INIT_1 = 16'h0000;
defparam ram16sdp_inst_143.INIT_2 = 16'h0000;
defparam ram16sdp_inst_143.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_144 (
    .DO(ram16sdp_inst_144_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_56),
    .CLK(clk)
);

defparam ram16sdp_inst_144.INIT_0 = 16'h0000;
defparam ram16sdp_inst_144.INIT_1 = 16'h0000;
defparam ram16sdp_inst_144.INIT_2 = 16'h0000;
defparam ram16sdp_inst_144.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_145 (
    .DO(ram16sdp_inst_145_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_56),
    .CLK(clk)
);

defparam ram16sdp_inst_145.INIT_0 = 16'h0000;
defparam ram16sdp_inst_145.INIT_1 = 16'h0000;
defparam ram16sdp_inst_145.INIT_2 = 16'h0000;
defparam ram16sdp_inst_145.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_146 (
    .DO(ram16sdp_inst_146_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_56),
    .CLK(clk)
);

defparam ram16sdp_inst_146.INIT_0 = 16'h0000;
defparam ram16sdp_inst_146.INIT_1 = 16'h0000;
defparam ram16sdp_inst_146.INIT_2 = 16'h0000;
defparam ram16sdp_inst_146.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_147 (
    .DO(ram16sdp_inst_147_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_56),
    .CLK(clk)
);

defparam ram16sdp_inst_147.INIT_0 = 16'h0000;
defparam ram16sdp_inst_147.INIT_1 = 16'h0000;
defparam ram16sdp_inst_147.INIT_2 = 16'h0000;
defparam ram16sdp_inst_147.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_148 (
    .DO(ram16sdp_inst_148_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_56),
    .CLK(clk)
);

defparam ram16sdp_inst_148.INIT_0 = 16'h0000;
defparam ram16sdp_inst_148.INIT_1 = 16'h0000;
defparam ram16sdp_inst_148.INIT_2 = 16'h0000;
defparam ram16sdp_inst_148.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_149 (
    .DO(ram16sdp_inst_149_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_56),
    .CLK(clk)
);

defparam ram16sdp_inst_149.INIT_0 = 16'h0000;
defparam ram16sdp_inst_149.INIT_1 = 16'h0000;
defparam ram16sdp_inst_149.INIT_2 = 16'h0000;
defparam ram16sdp_inst_149.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_150 (
    .DO(ram16sdp_inst_150_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_56),
    .CLK(clk)
);

defparam ram16sdp_inst_150.INIT_0 = 16'h0000;
defparam ram16sdp_inst_150.INIT_1 = 16'h0000;
defparam ram16sdp_inst_150.INIT_2 = 16'h0000;
defparam ram16sdp_inst_150.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_151 (
    .DO(ram16sdp_inst_151_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_56),
    .CLK(clk)
);

defparam ram16sdp_inst_151.INIT_0 = 16'h0000;
defparam ram16sdp_inst_151.INIT_1 = 16'h0000;
defparam ram16sdp_inst_151.INIT_2 = 16'h0000;
defparam ram16sdp_inst_151.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_152 (
    .DO(ram16sdp_inst_152_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_152.INIT_0 = 16'h0000;
defparam ram16sdp_inst_152.INIT_1 = 16'h0000;
defparam ram16sdp_inst_152.INIT_2 = 16'h0000;
defparam ram16sdp_inst_152.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_153 (
    .DO(ram16sdp_inst_153_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_153.INIT_0 = 16'h0000;
defparam ram16sdp_inst_153.INIT_1 = 16'h0000;
defparam ram16sdp_inst_153.INIT_2 = 16'h0000;
defparam ram16sdp_inst_153.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_154 (
    .DO(ram16sdp_inst_154_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_154.INIT_0 = 16'h0000;
defparam ram16sdp_inst_154.INIT_1 = 16'h0000;
defparam ram16sdp_inst_154.INIT_2 = 16'h0000;
defparam ram16sdp_inst_154.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_155 (
    .DO(ram16sdp_inst_155_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_155.INIT_0 = 16'h0000;
defparam ram16sdp_inst_155.INIT_1 = 16'h0000;
defparam ram16sdp_inst_155.INIT_2 = 16'h0000;
defparam ram16sdp_inst_155.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_156 (
    .DO(ram16sdp_inst_156_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_156.INIT_0 = 16'h0000;
defparam ram16sdp_inst_156.INIT_1 = 16'h0000;
defparam ram16sdp_inst_156.INIT_2 = 16'h0000;
defparam ram16sdp_inst_156.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_157 (
    .DO(ram16sdp_inst_157_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_157.INIT_0 = 16'h0000;
defparam ram16sdp_inst_157.INIT_1 = 16'h0000;
defparam ram16sdp_inst_157.INIT_2 = 16'h0000;
defparam ram16sdp_inst_157.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_158 (
    .DO(ram16sdp_inst_158_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_158.INIT_0 = 16'h0000;
defparam ram16sdp_inst_158.INIT_1 = 16'h0000;
defparam ram16sdp_inst_158.INIT_2 = 16'h0000;
defparam ram16sdp_inst_158.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_159 (
    .DO(ram16sdp_inst_159_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_159.INIT_0 = 16'h0000;
defparam ram16sdp_inst_159.INIT_1 = 16'h0000;
defparam ram16sdp_inst_159.INIT_2 = 16'h0000;
defparam ram16sdp_inst_159.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_160 (
    .DO(ram16sdp_inst_160_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_62),
    .CLK(clk)
);

defparam ram16sdp_inst_160.INIT_0 = 16'h0000;
defparam ram16sdp_inst_160.INIT_1 = 16'h0000;
defparam ram16sdp_inst_160.INIT_2 = 16'h0000;
defparam ram16sdp_inst_160.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_161 (
    .DO(ram16sdp_inst_161_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_62),
    .CLK(clk)
);

defparam ram16sdp_inst_161.INIT_0 = 16'h0000;
defparam ram16sdp_inst_161.INIT_1 = 16'h0000;
defparam ram16sdp_inst_161.INIT_2 = 16'h0000;
defparam ram16sdp_inst_161.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_162 (
    .DO(ram16sdp_inst_162_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_62),
    .CLK(clk)
);

defparam ram16sdp_inst_162.INIT_0 = 16'h0000;
defparam ram16sdp_inst_162.INIT_1 = 16'h0000;
defparam ram16sdp_inst_162.INIT_2 = 16'h0000;
defparam ram16sdp_inst_162.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_163 (
    .DO(ram16sdp_inst_163_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_62),
    .CLK(clk)
);

defparam ram16sdp_inst_163.INIT_0 = 16'h0000;
defparam ram16sdp_inst_163.INIT_1 = 16'h0000;
defparam ram16sdp_inst_163.INIT_2 = 16'h0000;
defparam ram16sdp_inst_163.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_164 (
    .DO(ram16sdp_inst_164_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_62),
    .CLK(clk)
);

defparam ram16sdp_inst_164.INIT_0 = 16'h0000;
defparam ram16sdp_inst_164.INIT_1 = 16'h0000;
defparam ram16sdp_inst_164.INIT_2 = 16'h0000;
defparam ram16sdp_inst_164.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_165 (
    .DO(ram16sdp_inst_165_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_62),
    .CLK(clk)
);

defparam ram16sdp_inst_165.INIT_0 = 16'h0000;
defparam ram16sdp_inst_165.INIT_1 = 16'h0000;
defparam ram16sdp_inst_165.INIT_2 = 16'h0000;
defparam ram16sdp_inst_165.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_166 (
    .DO(ram16sdp_inst_166_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_62),
    .CLK(clk)
);

defparam ram16sdp_inst_166.INIT_0 = 16'h0000;
defparam ram16sdp_inst_166.INIT_1 = 16'h0000;
defparam ram16sdp_inst_166.INIT_2 = 16'h0000;
defparam ram16sdp_inst_166.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_167 (
    .DO(ram16sdp_inst_167_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_62),
    .CLK(clk)
);

defparam ram16sdp_inst_167.INIT_0 = 16'h0000;
defparam ram16sdp_inst_167.INIT_1 = 16'h0000;
defparam ram16sdp_inst_167.INIT_2 = 16'h0000;
defparam ram16sdp_inst_167.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_168 (
    .DO(ram16sdp_inst_168_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_168.INIT_0 = 16'h0000;
defparam ram16sdp_inst_168.INIT_1 = 16'h0000;
defparam ram16sdp_inst_168.INIT_2 = 16'h0000;
defparam ram16sdp_inst_168.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_169 (
    .DO(ram16sdp_inst_169_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_169.INIT_0 = 16'h0000;
defparam ram16sdp_inst_169.INIT_1 = 16'h0000;
defparam ram16sdp_inst_169.INIT_2 = 16'h0000;
defparam ram16sdp_inst_169.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_170 (
    .DO(ram16sdp_inst_170_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_170.INIT_0 = 16'h0000;
defparam ram16sdp_inst_170.INIT_1 = 16'h0000;
defparam ram16sdp_inst_170.INIT_2 = 16'h0000;
defparam ram16sdp_inst_170.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_171 (
    .DO(ram16sdp_inst_171_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_171.INIT_0 = 16'h0000;
defparam ram16sdp_inst_171.INIT_1 = 16'h0000;
defparam ram16sdp_inst_171.INIT_2 = 16'h0000;
defparam ram16sdp_inst_171.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_172 (
    .DO(ram16sdp_inst_172_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_172.INIT_0 = 16'h0000;
defparam ram16sdp_inst_172.INIT_1 = 16'h0000;
defparam ram16sdp_inst_172.INIT_2 = 16'h0000;
defparam ram16sdp_inst_172.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_173 (
    .DO(ram16sdp_inst_173_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_173.INIT_0 = 16'h0000;
defparam ram16sdp_inst_173.INIT_1 = 16'h0000;
defparam ram16sdp_inst_173.INIT_2 = 16'h0000;
defparam ram16sdp_inst_173.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_174 (
    .DO(ram16sdp_inst_174_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_174.INIT_0 = 16'h0000;
defparam ram16sdp_inst_174.INIT_1 = 16'h0000;
defparam ram16sdp_inst_174.INIT_2 = 16'h0000;
defparam ram16sdp_inst_174.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_175 (
    .DO(ram16sdp_inst_175_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_175.INIT_0 = 16'h0000;
defparam ram16sdp_inst_175.INIT_1 = 16'h0000;
defparam ram16sdp_inst_175.INIT_2 = 16'h0000;
defparam ram16sdp_inst_175.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_176 (
    .DO(ram16sdp_inst_176_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_68),
    .CLK(clk)
);

defparam ram16sdp_inst_176.INIT_0 = 16'h0000;
defparam ram16sdp_inst_176.INIT_1 = 16'h0000;
defparam ram16sdp_inst_176.INIT_2 = 16'h0000;
defparam ram16sdp_inst_176.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_177 (
    .DO(ram16sdp_inst_177_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_68),
    .CLK(clk)
);

defparam ram16sdp_inst_177.INIT_0 = 16'h0000;
defparam ram16sdp_inst_177.INIT_1 = 16'h0000;
defparam ram16sdp_inst_177.INIT_2 = 16'h0000;
defparam ram16sdp_inst_177.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_178 (
    .DO(ram16sdp_inst_178_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_68),
    .CLK(clk)
);

defparam ram16sdp_inst_178.INIT_0 = 16'h0000;
defparam ram16sdp_inst_178.INIT_1 = 16'h0000;
defparam ram16sdp_inst_178.INIT_2 = 16'h0000;
defparam ram16sdp_inst_178.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_179 (
    .DO(ram16sdp_inst_179_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_68),
    .CLK(clk)
);

defparam ram16sdp_inst_179.INIT_0 = 16'h0000;
defparam ram16sdp_inst_179.INIT_1 = 16'h0000;
defparam ram16sdp_inst_179.INIT_2 = 16'h0000;
defparam ram16sdp_inst_179.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_180 (
    .DO(ram16sdp_inst_180_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_68),
    .CLK(clk)
);

defparam ram16sdp_inst_180.INIT_0 = 16'h0000;
defparam ram16sdp_inst_180.INIT_1 = 16'h0000;
defparam ram16sdp_inst_180.INIT_2 = 16'h0000;
defparam ram16sdp_inst_180.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_181 (
    .DO(ram16sdp_inst_181_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_68),
    .CLK(clk)
);

defparam ram16sdp_inst_181.INIT_0 = 16'h0000;
defparam ram16sdp_inst_181.INIT_1 = 16'h0000;
defparam ram16sdp_inst_181.INIT_2 = 16'h0000;
defparam ram16sdp_inst_181.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_182 (
    .DO(ram16sdp_inst_182_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_68),
    .CLK(clk)
);

defparam ram16sdp_inst_182.INIT_0 = 16'h0000;
defparam ram16sdp_inst_182.INIT_1 = 16'h0000;
defparam ram16sdp_inst_182.INIT_2 = 16'h0000;
defparam ram16sdp_inst_182.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_183 (
    .DO(ram16sdp_inst_183_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_68),
    .CLK(clk)
);

defparam ram16sdp_inst_183.INIT_0 = 16'h0000;
defparam ram16sdp_inst_183.INIT_1 = 16'h0000;
defparam ram16sdp_inst_183.INIT_2 = 16'h0000;
defparam ram16sdp_inst_183.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_184 (
    .DO(ram16sdp_inst_184_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_184.INIT_0 = 16'h0000;
defparam ram16sdp_inst_184.INIT_1 = 16'h0000;
defparam ram16sdp_inst_184.INIT_2 = 16'h0000;
defparam ram16sdp_inst_184.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_185 (
    .DO(ram16sdp_inst_185_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_185.INIT_0 = 16'h0000;
defparam ram16sdp_inst_185.INIT_1 = 16'h0000;
defparam ram16sdp_inst_185.INIT_2 = 16'h0000;
defparam ram16sdp_inst_185.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_186 (
    .DO(ram16sdp_inst_186_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_186.INIT_0 = 16'h0000;
defparam ram16sdp_inst_186.INIT_1 = 16'h0000;
defparam ram16sdp_inst_186.INIT_2 = 16'h0000;
defparam ram16sdp_inst_186.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_187 (
    .DO(ram16sdp_inst_187_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_187.INIT_0 = 16'h0000;
defparam ram16sdp_inst_187.INIT_1 = 16'h0000;
defparam ram16sdp_inst_187.INIT_2 = 16'h0000;
defparam ram16sdp_inst_187.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_188 (
    .DO(ram16sdp_inst_188_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_188.INIT_0 = 16'h0000;
defparam ram16sdp_inst_188.INIT_1 = 16'h0000;
defparam ram16sdp_inst_188.INIT_2 = 16'h0000;
defparam ram16sdp_inst_188.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_189 (
    .DO(ram16sdp_inst_189_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_189.INIT_0 = 16'h0000;
defparam ram16sdp_inst_189.INIT_1 = 16'h0000;
defparam ram16sdp_inst_189.INIT_2 = 16'h0000;
defparam ram16sdp_inst_189.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_190 (
    .DO(ram16sdp_inst_190_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_190.INIT_0 = 16'h0000;
defparam ram16sdp_inst_190.INIT_1 = 16'h0000;
defparam ram16sdp_inst_190.INIT_2 = 16'h0000;
defparam ram16sdp_inst_190.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_191 (
    .DO(ram16sdp_inst_191_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_191.INIT_0 = 16'h0000;
defparam ram16sdp_inst_191.INIT_1 = 16'h0000;
defparam ram16sdp_inst_191.INIT_2 = 16'h0000;
defparam ram16sdp_inst_191.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_192 (
    .DO(ram16sdp_inst_192_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_74),
    .CLK(clk)
);

defparam ram16sdp_inst_192.INIT_0 = 16'h0000;
defparam ram16sdp_inst_192.INIT_1 = 16'h0000;
defparam ram16sdp_inst_192.INIT_2 = 16'h0000;
defparam ram16sdp_inst_192.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_193 (
    .DO(ram16sdp_inst_193_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_74),
    .CLK(clk)
);

defparam ram16sdp_inst_193.INIT_0 = 16'h0000;
defparam ram16sdp_inst_193.INIT_1 = 16'h0000;
defparam ram16sdp_inst_193.INIT_2 = 16'h0000;
defparam ram16sdp_inst_193.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_194 (
    .DO(ram16sdp_inst_194_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_74),
    .CLK(clk)
);

defparam ram16sdp_inst_194.INIT_0 = 16'h0000;
defparam ram16sdp_inst_194.INIT_1 = 16'h0000;
defparam ram16sdp_inst_194.INIT_2 = 16'h0000;
defparam ram16sdp_inst_194.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_195 (
    .DO(ram16sdp_inst_195_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_74),
    .CLK(clk)
);

defparam ram16sdp_inst_195.INIT_0 = 16'h0000;
defparam ram16sdp_inst_195.INIT_1 = 16'h0000;
defparam ram16sdp_inst_195.INIT_2 = 16'h0000;
defparam ram16sdp_inst_195.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_196 (
    .DO(ram16sdp_inst_196_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_74),
    .CLK(clk)
);

defparam ram16sdp_inst_196.INIT_0 = 16'h0000;
defparam ram16sdp_inst_196.INIT_1 = 16'h0000;
defparam ram16sdp_inst_196.INIT_2 = 16'h0000;
defparam ram16sdp_inst_196.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_197 (
    .DO(ram16sdp_inst_197_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_74),
    .CLK(clk)
);

defparam ram16sdp_inst_197.INIT_0 = 16'h0000;
defparam ram16sdp_inst_197.INIT_1 = 16'h0000;
defparam ram16sdp_inst_197.INIT_2 = 16'h0000;
defparam ram16sdp_inst_197.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_198 (
    .DO(ram16sdp_inst_198_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_74),
    .CLK(clk)
);

defparam ram16sdp_inst_198.INIT_0 = 16'h0000;
defparam ram16sdp_inst_198.INIT_1 = 16'h0000;
defparam ram16sdp_inst_198.INIT_2 = 16'h0000;
defparam ram16sdp_inst_198.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_199 (
    .DO(ram16sdp_inst_199_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_74),
    .CLK(clk)
);

defparam ram16sdp_inst_199.INIT_0 = 16'h0000;
defparam ram16sdp_inst_199.INIT_1 = 16'h0000;
defparam ram16sdp_inst_199.INIT_2 = 16'h0000;
defparam ram16sdp_inst_199.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_200 (
    .DO(ram16sdp_inst_200_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_200.INIT_0 = 16'h0000;
defparam ram16sdp_inst_200.INIT_1 = 16'h0000;
defparam ram16sdp_inst_200.INIT_2 = 16'h0000;
defparam ram16sdp_inst_200.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_201 (
    .DO(ram16sdp_inst_201_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_201.INIT_0 = 16'h0000;
defparam ram16sdp_inst_201.INIT_1 = 16'h0000;
defparam ram16sdp_inst_201.INIT_2 = 16'h0000;
defparam ram16sdp_inst_201.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_202 (
    .DO(ram16sdp_inst_202_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_202.INIT_0 = 16'h0000;
defparam ram16sdp_inst_202.INIT_1 = 16'h0000;
defparam ram16sdp_inst_202.INIT_2 = 16'h0000;
defparam ram16sdp_inst_202.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_203 (
    .DO(ram16sdp_inst_203_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_203.INIT_0 = 16'h0000;
defparam ram16sdp_inst_203.INIT_1 = 16'h0000;
defparam ram16sdp_inst_203.INIT_2 = 16'h0000;
defparam ram16sdp_inst_203.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_204 (
    .DO(ram16sdp_inst_204_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_204.INIT_0 = 16'h0000;
defparam ram16sdp_inst_204.INIT_1 = 16'h0000;
defparam ram16sdp_inst_204.INIT_2 = 16'h0000;
defparam ram16sdp_inst_204.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_205 (
    .DO(ram16sdp_inst_205_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_205.INIT_0 = 16'h0000;
defparam ram16sdp_inst_205.INIT_1 = 16'h0000;
defparam ram16sdp_inst_205.INIT_2 = 16'h0000;
defparam ram16sdp_inst_205.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_206 (
    .DO(ram16sdp_inst_206_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_206.INIT_0 = 16'h0000;
defparam ram16sdp_inst_206.INIT_1 = 16'h0000;
defparam ram16sdp_inst_206.INIT_2 = 16'h0000;
defparam ram16sdp_inst_206.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_207 (
    .DO(ram16sdp_inst_207_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_207.INIT_0 = 16'h0000;
defparam ram16sdp_inst_207.INIT_1 = 16'h0000;
defparam ram16sdp_inst_207.INIT_2 = 16'h0000;
defparam ram16sdp_inst_207.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_208 (
    .DO(ram16sdp_inst_208_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_80),
    .CLK(clk)
);

defparam ram16sdp_inst_208.INIT_0 = 16'h0000;
defparam ram16sdp_inst_208.INIT_1 = 16'h0000;
defparam ram16sdp_inst_208.INIT_2 = 16'h0000;
defparam ram16sdp_inst_208.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_209 (
    .DO(ram16sdp_inst_209_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_80),
    .CLK(clk)
);

defparam ram16sdp_inst_209.INIT_0 = 16'h0000;
defparam ram16sdp_inst_209.INIT_1 = 16'h0000;
defparam ram16sdp_inst_209.INIT_2 = 16'h0000;
defparam ram16sdp_inst_209.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_210 (
    .DO(ram16sdp_inst_210_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_80),
    .CLK(clk)
);

defparam ram16sdp_inst_210.INIT_0 = 16'h0000;
defparam ram16sdp_inst_210.INIT_1 = 16'h0000;
defparam ram16sdp_inst_210.INIT_2 = 16'h0000;
defparam ram16sdp_inst_210.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_211 (
    .DO(ram16sdp_inst_211_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_80),
    .CLK(clk)
);

defparam ram16sdp_inst_211.INIT_0 = 16'h0000;
defparam ram16sdp_inst_211.INIT_1 = 16'h0000;
defparam ram16sdp_inst_211.INIT_2 = 16'h0000;
defparam ram16sdp_inst_211.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_212 (
    .DO(ram16sdp_inst_212_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_80),
    .CLK(clk)
);

defparam ram16sdp_inst_212.INIT_0 = 16'h0000;
defparam ram16sdp_inst_212.INIT_1 = 16'h0000;
defparam ram16sdp_inst_212.INIT_2 = 16'h0000;
defparam ram16sdp_inst_212.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_213 (
    .DO(ram16sdp_inst_213_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_80),
    .CLK(clk)
);

defparam ram16sdp_inst_213.INIT_0 = 16'h0000;
defparam ram16sdp_inst_213.INIT_1 = 16'h0000;
defparam ram16sdp_inst_213.INIT_2 = 16'h0000;
defparam ram16sdp_inst_213.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_214 (
    .DO(ram16sdp_inst_214_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_80),
    .CLK(clk)
);

defparam ram16sdp_inst_214.INIT_0 = 16'h0000;
defparam ram16sdp_inst_214.INIT_1 = 16'h0000;
defparam ram16sdp_inst_214.INIT_2 = 16'h0000;
defparam ram16sdp_inst_214.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_215 (
    .DO(ram16sdp_inst_215_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_80),
    .CLK(clk)
);

defparam ram16sdp_inst_215.INIT_0 = 16'h0000;
defparam ram16sdp_inst_215.INIT_1 = 16'h0000;
defparam ram16sdp_inst_215.INIT_2 = 16'h0000;
defparam ram16sdp_inst_215.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_216 (
    .DO(ram16sdp_inst_216_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_216.INIT_0 = 16'h0000;
defparam ram16sdp_inst_216.INIT_1 = 16'h0000;
defparam ram16sdp_inst_216.INIT_2 = 16'h0000;
defparam ram16sdp_inst_216.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_217 (
    .DO(ram16sdp_inst_217_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_217.INIT_0 = 16'h0000;
defparam ram16sdp_inst_217.INIT_1 = 16'h0000;
defparam ram16sdp_inst_217.INIT_2 = 16'h0000;
defparam ram16sdp_inst_217.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_218 (
    .DO(ram16sdp_inst_218_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_218.INIT_0 = 16'h0000;
defparam ram16sdp_inst_218.INIT_1 = 16'h0000;
defparam ram16sdp_inst_218.INIT_2 = 16'h0000;
defparam ram16sdp_inst_218.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_219 (
    .DO(ram16sdp_inst_219_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_219.INIT_0 = 16'h0000;
defparam ram16sdp_inst_219.INIT_1 = 16'h0000;
defparam ram16sdp_inst_219.INIT_2 = 16'h0000;
defparam ram16sdp_inst_219.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_220 (
    .DO(ram16sdp_inst_220_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_220.INIT_0 = 16'h0000;
defparam ram16sdp_inst_220.INIT_1 = 16'h0000;
defparam ram16sdp_inst_220.INIT_2 = 16'h0000;
defparam ram16sdp_inst_220.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_221 (
    .DO(ram16sdp_inst_221_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_221.INIT_0 = 16'h0000;
defparam ram16sdp_inst_221.INIT_1 = 16'h0000;
defparam ram16sdp_inst_221.INIT_2 = 16'h0000;
defparam ram16sdp_inst_221.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_222 (
    .DO(ram16sdp_inst_222_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_222.INIT_0 = 16'h0000;
defparam ram16sdp_inst_222.INIT_1 = 16'h0000;
defparam ram16sdp_inst_222.INIT_2 = 16'h0000;
defparam ram16sdp_inst_222.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_223 (
    .DO(ram16sdp_inst_223_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_223.INIT_0 = 16'h0000;
defparam ram16sdp_inst_223.INIT_1 = 16'h0000;
defparam ram16sdp_inst_223.INIT_2 = 16'h0000;
defparam ram16sdp_inst_223.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_224 (
    .DO(ram16sdp_inst_224_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_86),
    .CLK(clk)
);

defparam ram16sdp_inst_224.INIT_0 = 16'h0000;
defparam ram16sdp_inst_224.INIT_1 = 16'h0000;
defparam ram16sdp_inst_224.INIT_2 = 16'h0000;
defparam ram16sdp_inst_224.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_225 (
    .DO(ram16sdp_inst_225_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_86),
    .CLK(clk)
);

defparam ram16sdp_inst_225.INIT_0 = 16'h0000;
defparam ram16sdp_inst_225.INIT_1 = 16'h0000;
defparam ram16sdp_inst_225.INIT_2 = 16'h0000;
defparam ram16sdp_inst_225.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_226 (
    .DO(ram16sdp_inst_226_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_86),
    .CLK(clk)
);

defparam ram16sdp_inst_226.INIT_0 = 16'h0000;
defparam ram16sdp_inst_226.INIT_1 = 16'h0000;
defparam ram16sdp_inst_226.INIT_2 = 16'h0000;
defparam ram16sdp_inst_226.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_227 (
    .DO(ram16sdp_inst_227_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_86),
    .CLK(clk)
);

defparam ram16sdp_inst_227.INIT_0 = 16'h0000;
defparam ram16sdp_inst_227.INIT_1 = 16'h0000;
defparam ram16sdp_inst_227.INIT_2 = 16'h0000;
defparam ram16sdp_inst_227.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_228 (
    .DO(ram16sdp_inst_228_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_86),
    .CLK(clk)
);

defparam ram16sdp_inst_228.INIT_0 = 16'h0000;
defparam ram16sdp_inst_228.INIT_1 = 16'h0000;
defparam ram16sdp_inst_228.INIT_2 = 16'h0000;
defparam ram16sdp_inst_228.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_229 (
    .DO(ram16sdp_inst_229_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_86),
    .CLK(clk)
);

defparam ram16sdp_inst_229.INIT_0 = 16'h0000;
defparam ram16sdp_inst_229.INIT_1 = 16'h0000;
defparam ram16sdp_inst_229.INIT_2 = 16'h0000;
defparam ram16sdp_inst_229.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_230 (
    .DO(ram16sdp_inst_230_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_86),
    .CLK(clk)
);

defparam ram16sdp_inst_230.INIT_0 = 16'h0000;
defparam ram16sdp_inst_230.INIT_1 = 16'h0000;
defparam ram16sdp_inst_230.INIT_2 = 16'h0000;
defparam ram16sdp_inst_230.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_231 (
    .DO(ram16sdp_inst_231_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_86),
    .CLK(clk)
);

defparam ram16sdp_inst_231.INIT_0 = 16'h0000;
defparam ram16sdp_inst_231.INIT_1 = 16'h0000;
defparam ram16sdp_inst_231.INIT_2 = 16'h0000;
defparam ram16sdp_inst_231.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_232 (
    .DO(ram16sdp_inst_232_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_232.INIT_0 = 16'h0000;
defparam ram16sdp_inst_232.INIT_1 = 16'h0000;
defparam ram16sdp_inst_232.INIT_2 = 16'h0000;
defparam ram16sdp_inst_232.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_233 (
    .DO(ram16sdp_inst_233_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_233.INIT_0 = 16'h0000;
defparam ram16sdp_inst_233.INIT_1 = 16'h0000;
defparam ram16sdp_inst_233.INIT_2 = 16'h0000;
defparam ram16sdp_inst_233.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_234 (
    .DO(ram16sdp_inst_234_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_234.INIT_0 = 16'h0000;
defparam ram16sdp_inst_234.INIT_1 = 16'h0000;
defparam ram16sdp_inst_234.INIT_2 = 16'h0000;
defparam ram16sdp_inst_234.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_235 (
    .DO(ram16sdp_inst_235_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_235.INIT_0 = 16'h0000;
defparam ram16sdp_inst_235.INIT_1 = 16'h0000;
defparam ram16sdp_inst_235.INIT_2 = 16'h0000;
defparam ram16sdp_inst_235.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_236 (
    .DO(ram16sdp_inst_236_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_236.INIT_0 = 16'h0000;
defparam ram16sdp_inst_236.INIT_1 = 16'h0000;
defparam ram16sdp_inst_236.INIT_2 = 16'h0000;
defparam ram16sdp_inst_236.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_237 (
    .DO(ram16sdp_inst_237_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_237.INIT_0 = 16'h0000;
defparam ram16sdp_inst_237.INIT_1 = 16'h0000;
defparam ram16sdp_inst_237.INIT_2 = 16'h0000;
defparam ram16sdp_inst_237.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_238 (
    .DO(ram16sdp_inst_238_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_238.INIT_0 = 16'h0000;
defparam ram16sdp_inst_238.INIT_1 = 16'h0000;
defparam ram16sdp_inst_238.INIT_2 = 16'h0000;
defparam ram16sdp_inst_238.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_239 (
    .DO(ram16sdp_inst_239_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_239.INIT_0 = 16'h0000;
defparam ram16sdp_inst_239.INIT_1 = 16'h0000;
defparam ram16sdp_inst_239.INIT_2 = 16'h0000;
defparam ram16sdp_inst_239.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_240 (
    .DO(ram16sdp_inst_240_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_92),
    .CLK(clk)
);

defparam ram16sdp_inst_240.INIT_0 = 16'h0000;
defparam ram16sdp_inst_240.INIT_1 = 16'h0000;
defparam ram16sdp_inst_240.INIT_2 = 16'h0000;
defparam ram16sdp_inst_240.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_241 (
    .DO(ram16sdp_inst_241_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_92),
    .CLK(clk)
);

defparam ram16sdp_inst_241.INIT_0 = 16'h0000;
defparam ram16sdp_inst_241.INIT_1 = 16'h0000;
defparam ram16sdp_inst_241.INIT_2 = 16'h0000;
defparam ram16sdp_inst_241.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_242 (
    .DO(ram16sdp_inst_242_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_92),
    .CLK(clk)
);

defparam ram16sdp_inst_242.INIT_0 = 16'h0000;
defparam ram16sdp_inst_242.INIT_1 = 16'h0000;
defparam ram16sdp_inst_242.INIT_2 = 16'h0000;
defparam ram16sdp_inst_242.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_243 (
    .DO(ram16sdp_inst_243_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_92),
    .CLK(clk)
);

defparam ram16sdp_inst_243.INIT_0 = 16'h0000;
defparam ram16sdp_inst_243.INIT_1 = 16'h0000;
defparam ram16sdp_inst_243.INIT_2 = 16'h0000;
defparam ram16sdp_inst_243.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_244 (
    .DO(ram16sdp_inst_244_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_92),
    .CLK(clk)
);

defparam ram16sdp_inst_244.INIT_0 = 16'h0000;
defparam ram16sdp_inst_244.INIT_1 = 16'h0000;
defparam ram16sdp_inst_244.INIT_2 = 16'h0000;
defparam ram16sdp_inst_244.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_245 (
    .DO(ram16sdp_inst_245_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_92),
    .CLK(clk)
);

defparam ram16sdp_inst_245.INIT_0 = 16'h0000;
defparam ram16sdp_inst_245.INIT_1 = 16'h0000;
defparam ram16sdp_inst_245.INIT_2 = 16'h0000;
defparam ram16sdp_inst_245.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_246 (
    .DO(ram16sdp_inst_246_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_92),
    .CLK(clk)
);

defparam ram16sdp_inst_246.INIT_0 = 16'h0000;
defparam ram16sdp_inst_246.INIT_1 = 16'h0000;
defparam ram16sdp_inst_246.INIT_2 = 16'h0000;
defparam ram16sdp_inst_246.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_247 (
    .DO(ram16sdp_inst_247_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_92),
    .CLK(clk)
);

defparam ram16sdp_inst_247.INIT_0 = 16'h0000;
defparam ram16sdp_inst_247.INIT_1 = 16'h0000;
defparam ram16sdp_inst_247.INIT_2 = 16'h0000;
defparam ram16sdp_inst_247.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_248 (
    .DO(ram16sdp_inst_248_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_248.INIT_0 = 16'h0000;
defparam ram16sdp_inst_248.INIT_1 = 16'h0000;
defparam ram16sdp_inst_248.INIT_2 = 16'h0000;
defparam ram16sdp_inst_248.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_249 (
    .DO(ram16sdp_inst_249_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_249.INIT_0 = 16'h0000;
defparam ram16sdp_inst_249.INIT_1 = 16'h0000;
defparam ram16sdp_inst_249.INIT_2 = 16'h0000;
defparam ram16sdp_inst_249.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_250 (
    .DO(ram16sdp_inst_250_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_250.INIT_0 = 16'h0000;
defparam ram16sdp_inst_250.INIT_1 = 16'h0000;
defparam ram16sdp_inst_250.INIT_2 = 16'h0000;
defparam ram16sdp_inst_250.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_251 (
    .DO(ram16sdp_inst_251_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_251.INIT_0 = 16'h0000;
defparam ram16sdp_inst_251.INIT_1 = 16'h0000;
defparam ram16sdp_inst_251.INIT_2 = 16'h0000;
defparam ram16sdp_inst_251.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_252 (
    .DO(ram16sdp_inst_252_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_252.INIT_0 = 16'h0000;
defparam ram16sdp_inst_252.INIT_1 = 16'h0000;
defparam ram16sdp_inst_252.INIT_2 = 16'h0000;
defparam ram16sdp_inst_252.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_253 (
    .DO(ram16sdp_inst_253_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_253.INIT_0 = 16'h0000;
defparam ram16sdp_inst_253.INIT_1 = 16'h0000;
defparam ram16sdp_inst_253.INIT_2 = 16'h0000;
defparam ram16sdp_inst_253.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_254 (
    .DO(ram16sdp_inst_254_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_254.INIT_0 = 16'h0000;
defparam ram16sdp_inst_254.INIT_1 = 16'h0000;
defparam ram16sdp_inst_254.INIT_2 = 16'h0000;
defparam ram16sdp_inst_254.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_255 (
    .DO(ram16sdp_inst_255_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_255.INIT_0 = 16'h0000;
defparam ram16sdp_inst_255.INIT_1 = 16'h0000;
defparam ram16sdp_inst_255.INIT_2 = 16'h0000;
defparam ram16sdp_inst_255.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_256 (
    .DO(ram16sdp_inst_256_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_98),
    .CLK(clk)
);

defparam ram16sdp_inst_256.INIT_0 = 16'h0000;
defparam ram16sdp_inst_256.INIT_1 = 16'h0000;
defparam ram16sdp_inst_256.INIT_2 = 16'h0000;
defparam ram16sdp_inst_256.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_257 (
    .DO(ram16sdp_inst_257_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_98),
    .CLK(clk)
);

defparam ram16sdp_inst_257.INIT_0 = 16'h0000;
defparam ram16sdp_inst_257.INIT_1 = 16'h0000;
defparam ram16sdp_inst_257.INIT_2 = 16'h0000;
defparam ram16sdp_inst_257.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_258 (
    .DO(ram16sdp_inst_258_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_98),
    .CLK(clk)
);

defparam ram16sdp_inst_258.INIT_0 = 16'h0000;
defparam ram16sdp_inst_258.INIT_1 = 16'h0000;
defparam ram16sdp_inst_258.INIT_2 = 16'h0000;
defparam ram16sdp_inst_258.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_259 (
    .DO(ram16sdp_inst_259_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_98),
    .CLK(clk)
);

defparam ram16sdp_inst_259.INIT_0 = 16'h0000;
defparam ram16sdp_inst_259.INIT_1 = 16'h0000;
defparam ram16sdp_inst_259.INIT_2 = 16'h0000;
defparam ram16sdp_inst_259.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_260 (
    .DO(ram16sdp_inst_260_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_98),
    .CLK(clk)
);

defparam ram16sdp_inst_260.INIT_0 = 16'h0000;
defparam ram16sdp_inst_260.INIT_1 = 16'h0000;
defparam ram16sdp_inst_260.INIT_2 = 16'h0000;
defparam ram16sdp_inst_260.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_261 (
    .DO(ram16sdp_inst_261_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_98),
    .CLK(clk)
);

defparam ram16sdp_inst_261.INIT_0 = 16'h0000;
defparam ram16sdp_inst_261.INIT_1 = 16'h0000;
defparam ram16sdp_inst_261.INIT_2 = 16'h0000;
defparam ram16sdp_inst_261.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_262 (
    .DO(ram16sdp_inst_262_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_98),
    .CLK(clk)
);

defparam ram16sdp_inst_262.INIT_0 = 16'h0000;
defparam ram16sdp_inst_262.INIT_1 = 16'h0000;
defparam ram16sdp_inst_262.INIT_2 = 16'h0000;
defparam ram16sdp_inst_262.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_263 (
    .DO(ram16sdp_inst_263_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_98),
    .CLK(clk)
);

defparam ram16sdp_inst_263.INIT_0 = 16'h0000;
defparam ram16sdp_inst_263.INIT_1 = 16'h0000;
defparam ram16sdp_inst_263.INIT_2 = 16'h0000;
defparam ram16sdp_inst_263.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_264 (
    .DO(ram16sdp_inst_264_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_101),
    .CLK(clk)
);

defparam ram16sdp_inst_264.INIT_0 = 16'h0000;
defparam ram16sdp_inst_264.INIT_1 = 16'h0000;
defparam ram16sdp_inst_264.INIT_2 = 16'h0000;
defparam ram16sdp_inst_264.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_265 (
    .DO(ram16sdp_inst_265_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_101),
    .CLK(clk)
);

defparam ram16sdp_inst_265.INIT_0 = 16'h0000;
defparam ram16sdp_inst_265.INIT_1 = 16'h0000;
defparam ram16sdp_inst_265.INIT_2 = 16'h0000;
defparam ram16sdp_inst_265.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_266 (
    .DO(ram16sdp_inst_266_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_101),
    .CLK(clk)
);

defparam ram16sdp_inst_266.INIT_0 = 16'h0000;
defparam ram16sdp_inst_266.INIT_1 = 16'h0000;
defparam ram16sdp_inst_266.INIT_2 = 16'h0000;
defparam ram16sdp_inst_266.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_267 (
    .DO(ram16sdp_inst_267_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_101),
    .CLK(clk)
);

defparam ram16sdp_inst_267.INIT_0 = 16'h0000;
defparam ram16sdp_inst_267.INIT_1 = 16'h0000;
defparam ram16sdp_inst_267.INIT_2 = 16'h0000;
defparam ram16sdp_inst_267.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_268 (
    .DO(ram16sdp_inst_268_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_101),
    .CLK(clk)
);

defparam ram16sdp_inst_268.INIT_0 = 16'h0000;
defparam ram16sdp_inst_268.INIT_1 = 16'h0000;
defparam ram16sdp_inst_268.INIT_2 = 16'h0000;
defparam ram16sdp_inst_268.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_269 (
    .DO(ram16sdp_inst_269_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_101),
    .CLK(clk)
);

defparam ram16sdp_inst_269.INIT_0 = 16'h0000;
defparam ram16sdp_inst_269.INIT_1 = 16'h0000;
defparam ram16sdp_inst_269.INIT_2 = 16'h0000;
defparam ram16sdp_inst_269.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_270 (
    .DO(ram16sdp_inst_270_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_101),
    .CLK(clk)
);

defparam ram16sdp_inst_270.INIT_0 = 16'h0000;
defparam ram16sdp_inst_270.INIT_1 = 16'h0000;
defparam ram16sdp_inst_270.INIT_2 = 16'h0000;
defparam ram16sdp_inst_270.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_271 (
    .DO(ram16sdp_inst_271_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_101),
    .CLK(clk)
);

defparam ram16sdp_inst_271.INIT_0 = 16'h0000;
defparam ram16sdp_inst_271.INIT_1 = 16'h0000;
defparam ram16sdp_inst_271.INIT_2 = 16'h0000;
defparam ram16sdp_inst_271.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_272 (
    .DO(ram16sdp_inst_272_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_104),
    .CLK(clk)
);

defparam ram16sdp_inst_272.INIT_0 = 16'h0000;
defparam ram16sdp_inst_272.INIT_1 = 16'h0000;
defparam ram16sdp_inst_272.INIT_2 = 16'h0000;
defparam ram16sdp_inst_272.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_273 (
    .DO(ram16sdp_inst_273_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_104),
    .CLK(clk)
);

defparam ram16sdp_inst_273.INIT_0 = 16'h0000;
defparam ram16sdp_inst_273.INIT_1 = 16'h0000;
defparam ram16sdp_inst_273.INIT_2 = 16'h0000;
defparam ram16sdp_inst_273.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_274 (
    .DO(ram16sdp_inst_274_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_104),
    .CLK(clk)
);

defparam ram16sdp_inst_274.INIT_0 = 16'h0000;
defparam ram16sdp_inst_274.INIT_1 = 16'h0000;
defparam ram16sdp_inst_274.INIT_2 = 16'h0000;
defparam ram16sdp_inst_274.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_275 (
    .DO(ram16sdp_inst_275_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_104),
    .CLK(clk)
);

defparam ram16sdp_inst_275.INIT_0 = 16'h0000;
defparam ram16sdp_inst_275.INIT_1 = 16'h0000;
defparam ram16sdp_inst_275.INIT_2 = 16'h0000;
defparam ram16sdp_inst_275.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_276 (
    .DO(ram16sdp_inst_276_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_104),
    .CLK(clk)
);

defparam ram16sdp_inst_276.INIT_0 = 16'h0000;
defparam ram16sdp_inst_276.INIT_1 = 16'h0000;
defparam ram16sdp_inst_276.INIT_2 = 16'h0000;
defparam ram16sdp_inst_276.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_277 (
    .DO(ram16sdp_inst_277_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_104),
    .CLK(clk)
);

defparam ram16sdp_inst_277.INIT_0 = 16'h0000;
defparam ram16sdp_inst_277.INIT_1 = 16'h0000;
defparam ram16sdp_inst_277.INIT_2 = 16'h0000;
defparam ram16sdp_inst_277.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_278 (
    .DO(ram16sdp_inst_278_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_104),
    .CLK(clk)
);

defparam ram16sdp_inst_278.INIT_0 = 16'h0000;
defparam ram16sdp_inst_278.INIT_1 = 16'h0000;
defparam ram16sdp_inst_278.INIT_2 = 16'h0000;
defparam ram16sdp_inst_278.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_279 (
    .DO(ram16sdp_inst_279_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_104),
    .CLK(clk)
);

defparam ram16sdp_inst_279.INIT_0 = 16'h0000;
defparam ram16sdp_inst_279.INIT_1 = 16'h0000;
defparam ram16sdp_inst_279.INIT_2 = 16'h0000;
defparam ram16sdp_inst_279.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_280 (
    .DO(ram16sdp_inst_280_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16sdp_inst_280.INIT_0 = 16'h0000;
defparam ram16sdp_inst_280.INIT_1 = 16'h0000;
defparam ram16sdp_inst_280.INIT_2 = 16'h0000;
defparam ram16sdp_inst_280.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_281 (
    .DO(ram16sdp_inst_281_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16sdp_inst_281.INIT_0 = 16'h0000;
defparam ram16sdp_inst_281.INIT_1 = 16'h0000;
defparam ram16sdp_inst_281.INIT_2 = 16'h0000;
defparam ram16sdp_inst_281.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_282 (
    .DO(ram16sdp_inst_282_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16sdp_inst_282.INIT_0 = 16'h0000;
defparam ram16sdp_inst_282.INIT_1 = 16'h0000;
defparam ram16sdp_inst_282.INIT_2 = 16'h0000;
defparam ram16sdp_inst_282.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_283 (
    .DO(ram16sdp_inst_283_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16sdp_inst_283.INIT_0 = 16'h0000;
defparam ram16sdp_inst_283.INIT_1 = 16'h0000;
defparam ram16sdp_inst_283.INIT_2 = 16'h0000;
defparam ram16sdp_inst_283.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_284 (
    .DO(ram16sdp_inst_284_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16sdp_inst_284.INIT_0 = 16'h0000;
defparam ram16sdp_inst_284.INIT_1 = 16'h0000;
defparam ram16sdp_inst_284.INIT_2 = 16'h0000;
defparam ram16sdp_inst_284.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_285 (
    .DO(ram16sdp_inst_285_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16sdp_inst_285.INIT_0 = 16'h0000;
defparam ram16sdp_inst_285.INIT_1 = 16'h0000;
defparam ram16sdp_inst_285.INIT_2 = 16'h0000;
defparam ram16sdp_inst_285.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_286 (
    .DO(ram16sdp_inst_286_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16sdp_inst_286.INIT_0 = 16'h0000;
defparam ram16sdp_inst_286.INIT_1 = 16'h0000;
defparam ram16sdp_inst_286.INIT_2 = 16'h0000;
defparam ram16sdp_inst_286.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_287 (
    .DO(ram16sdp_inst_287_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16sdp_inst_287.INIT_0 = 16'h0000;
defparam ram16sdp_inst_287.INIT_1 = 16'h0000;
defparam ram16sdp_inst_287.INIT_2 = 16'h0000;
defparam ram16sdp_inst_287.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_288 (
    .DO(ram16sdp_inst_288_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_110),
    .CLK(clk)
);

defparam ram16sdp_inst_288.INIT_0 = 16'h0000;
defparam ram16sdp_inst_288.INIT_1 = 16'h0000;
defparam ram16sdp_inst_288.INIT_2 = 16'h0000;
defparam ram16sdp_inst_288.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_289 (
    .DO(ram16sdp_inst_289_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_110),
    .CLK(clk)
);

defparam ram16sdp_inst_289.INIT_0 = 16'h0000;
defparam ram16sdp_inst_289.INIT_1 = 16'h0000;
defparam ram16sdp_inst_289.INIT_2 = 16'h0000;
defparam ram16sdp_inst_289.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_290 (
    .DO(ram16sdp_inst_290_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_110),
    .CLK(clk)
);

defparam ram16sdp_inst_290.INIT_0 = 16'h0000;
defparam ram16sdp_inst_290.INIT_1 = 16'h0000;
defparam ram16sdp_inst_290.INIT_2 = 16'h0000;
defparam ram16sdp_inst_290.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_291 (
    .DO(ram16sdp_inst_291_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_110),
    .CLK(clk)
);

defparam ram16sdp_inst_291.INIT_0 = 16'h0000;
defparam ram16sdp_inst_291.INIT_1 = 16'h0000;
defparam ram16sdp_inst_291.INIT_2 = 16'h0000;
defparam ram16sdp_inst_291.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_292 (
    .DO(ram16sdp_inst_292_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_110),
    .CLK(clk)
);

defparam ram16sdp_inst_292.INIT_0 = 16'h0000;
defparam ram16sdp_inst_292.INIT_1 = 16'h0000;
defparam ram16sdp_inst_292.INIT_2 = 16'h0000;
defparam ram16sdp_inst_292.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_293 (
    .DO(ram16sdp_inst_293_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_110),
    .CLK(clk)
);

defparam ram16sdp_inst_293.INIT_0 = 16'h0000;
defparam ram16sdp_inst_293.INIT_1 = 16'h0000;
defparam ram16sdp_inst_293.INIT_2 = 16'h0000;
defparam ram16sdp_inst_293.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_294 (
    .DO(ram16sdp_inst_294_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_110),
    .CLK(clk)
);

defparam ram16sdp_inst_294.INIT_0 = 16'h0000;
defparam ram16sdp_inst_294.INIT_1 = 16'h0000;
defparam ram16sdp_inst_294.INIT_2 = 16'h0000;
defparam ram16sdp_inst_294.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_295 (
    .DO(ram16sdp_inst_295_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_110),
    .CLK(clk)
);

defparam ram16sdp_inst_295.INIT_0 = 16'h0000;
defparam ram16sdp_inst_295.INIT_1 = 16'h0000;
defparam ram16sdp_inst_295.INIT_2 = 16'h0000;
defparam ram16sdp_inst_295.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_296 (
    .DO(ram16sdp_inst_296_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_113),
    .CLK(clk)
);

defparam ram16sdp_inst_296.INIT_0 = 16'h0000;
defparam ram16sdp_inst_296.INIT_1 = 16'h0000;
defparam ram16sdp_inst_296.INIT_2 = 16'h0000;
defparam ram16sdp_inst_296.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_297 (
    .DO(ram16sdp_inst_297_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_113),
    .CLK(clk)
);

defparam ram16sdp_inst_297.INIT_0 = 16'h0000;
defparam ram16sdp_inst_297.INIT_1 = 16'h0000;
defparam ram16sdp_inst_297.INIT_2 = 16'h0000;
defparam ram16sdp_inst_297.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_298 (
    .DO(ram16sdp_inst_298_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_113),
    .CLK(clk)
);

defparam ram16sdp_inst_298.INIT_0 = 16'h0000;
defparam ram16sdp_inst_298.INIT_1 = 16'h0000;
defparam ram16sdp_inst_298.INIT_2 = 16'h0000;
defparam ram16sdp_inst_298.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_299 (
    .DO(ram16sdp_inst_299_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_113),
    .CLK(clk)
);

defparam ram16sdp_inst_299.INIT_0 = 16'h0000;
defparam ram16sdp_inst_299.INIT_1 = 16'h0000;
defparam ram16sdp_inst_299.INIT_2 = 16'h0000;
defparam ram16sdp_inst_299.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_300 (
    .DO(ram16sdp_inst_300_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_113),
    .CLK(clk)
);

defparam ram16sdp_inst_300.INIT_0 = 16'h0000;
defparam ram16sdp_inst_300.INIT_1 = 16'h0000;
defparam ram16sdp_inst_300.INIT_2 = 16'h0000;
defparam ram16sdp_inst_300.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_301 (
    .DO(ram16sdp_inst_301_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_113),
    .CLK(clk)
);

defparam ram16sdp_inst_301.INIT_0 = 16'h0000;
defparam ram16sdp_inst_301.INIT_1 = 16'h0000;
defparam ram16sdp_inst_301.INIT_2 = 16'h0000;
defparam ram16sdp_inst_301.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_302 (
    .DO(ram16sdp_inst_302_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_113),
    .CLK(clk)
);

defparam ram16sdp_inst_302.INIT_0 = 16'h0000;
defparam ram16sdp_inst_302.INIT_1 = 16'h0000;
defparam ram16sdp_inst_302.INIT_2 = 16'h0000;
defparam ram16sdp_inst_302.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_303 (
    .DO(ram16sdp_inst_303_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_113),
    .CLK(clk)
);

defparam ram16sdp_inst_303.INIT_0 = 16'h0000;
defparam ram16sdp_inst_303.INIT_1 = 16'h0000;
defparam ram16sdp_inst_303.INIT_2 = 16'h0000;
defparam ram16sdp_inst_303.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_304 (
    .DO(ram16sdp_inst_304_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_116),
    .CLK(clk)
);

defparam ram16sdp_inst_304.INIT_0 = 16'h0000;
defparam ram16sdp_inst_304.INIT_1 = 16'h0000;
defparam ram16sdp_inst_304.INIT_2 = 16'h0000;
defparam ram16sdp_inst_304.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_305 (
    .DO(ram16sdp_inst_305_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_116),
    .CLK(clk)
);

defparam ram16sdp_inst_305.INIT_0 = 16'h0000;
defparam ram16sdp_inst_305.INIT_1 = 16'h0000;
defparam ram16sdp_inst_305.INIT_2 = 16'h0000;
defparam ram16sdp_inst_305.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_306 (
    .DO(ram16sdp_inst_306_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_116),
    .CLK(clk)
);

defparam ram16sdp_inst_306.INIT_0 = 16'h0000;
defparam ram16sdp_inst_306.INIT_1 = 16'h0000;
defparam ram16sdp_inst_306.INIT_2 = 16'h0000;
defparam ram16sdp_inst_306.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_307 (
    .DO(ram16sdp_inst_307_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_116),
    .CLK(clk)
);

defparam ram16sdp_inst_307.INIT_0 = 16'h0000;
defparam ram16sdp_inst_307.INIT_1 = 16'h0000;
defparam ram16sdp_inst_307.INIT_2 = 16'h0000;
defparam ram16sdp_inst_307.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_308 (
    .DO(ram16sdp_inst_308_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_116),
    .CLK(clk)
);

defparam ram16sdp_inst_308.INIT_0 = 16'h0000;
defparam ram16sdp_inst_308.INIT_1 = 16'h0000;
defparam ram16sdp_inst_308.INIT_2 = 16'h0000;
defparam ram16sdp_inst_308.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_309 (
    .DO(ram16sdp_inst_309_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_116),
    .CLK(clk)
);

defparam ram16sdp_inst_309.INIT_0 = 16'h0000;
defparam ram16sdp_inst_309.INIT_1 = 16'h0000;
defparam ram16sdp_inst_309.INIT_2 = 16'h0000;
defparam ram16sdp_inst_309.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_310 (
    .DO(ram16sdp_inst_310_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_116),
    .CLK(clk)
);

defparam ram16sdp_inst_310.INIT_0 = 16'h0000;
defparam ram16sdp_inst_310.INIT_1 = 16'h0000;
defparam ram16sdp_inst_310.INIT_2 = 16'h0000;
defparam ram16sdp_inst_310.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_311 (
    .DO(ram16sdp_inst_311_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_116),
    .CLK(clk)
);

defparam ram16sdp_inst_311.INIT_0 = 16'h0000;
defparam ram16sdp_inst_311.INIT_1 = 16'h0000;
defparam ram16sdp_inst_311.INIT_2 = 16'h0000;
defparam ram16sdp_inst_311.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_312 (
    .DO(ram16sdp_inst_312_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16sdp_inst_312.INIT_0 = 16'h0000;
defparam ram16sdp_inst_312.INIT_1 = 16'h0000;
defparam ram16sdp_inst_312.INIT_2 = 16'h0000;
defparam ram16sdp_inst_312.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_313 (
    .DO(ram16sdp_inst_313_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16sdp_inst_313.INIT_0 = 16'h0000;
defparam ram16sdp_inst_313.INIT_1 = 16'h0000;
defparam ram16sdp_inst_313.INIT_2 = 16'h0000;
defparam ram16sdp_inst_313.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_314 (
    .DO(ram16sdp_inst_314_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16sdp_inst_314.INIT_0 = 16'h0000;
defparam ram16sdp_inst_314.INIT_1 = 16'h0000;
defparam ram16sdp_inst_314.INIT_2 = 16'h0000;
defparam ram16sdp_inst_314.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_315 (
    .DO(ram16sdp_inst_315_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16sdp_inst_315.INIT_0 = 16'h0000;
defparam ram16sdp_inst_315.INIT_1 = 16'h0000;
defparam ram16sdp_inst_315.INIT_2 = 16'h0000;
defparam ram16sdp_inst_315.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_316 (
    .DO(ram16sdp_inst_316_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16sdp_inst_316.INIT_0 = 16'h0000;
defparam ram16sdp_inst_316.INIT_1 = 16'h0000;
defparam ram16sdp_inst_316.INIT_2 = 16'h0000;
defparam ram16sdp_inst_316.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_317 (
    .DO(ram16sdp_inst_317_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16sdp_inst_317.INIT_0 = 16'h0000;
defparam ram16sdp_inst_317.INIT_1 = 16'h0000;
defparam ram16sdp_inst_317.INIT_2 = 16'h0000;
defparam ram16sdp_inst_317.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_318 (
    .DO(ram16sdp_inst_318_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16sdp_inst_318.INIT_0 = 16'h0000;
defparam ram16sdp_inst_318.INIT_1 = 16'h0000;
defparam ram16sdp_inst_318.INIT_2 = 16'h0000;
defparam ram16sdp_inst_318.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_319 (
    .DO(ram16sdp_inst_319_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16sdp_inst_319.INIT_0 = 16'h0000;
defparam ram16sdp_inst_319.INIT_1 = 16'h0000;
defparam ram16sdp_inst_319.INIT_2 = 16'h0000;
defparam ram16sdp_inst_319.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_320 (
    .DO(ram16sdp_inst_320_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_122),
    .CLK(clk)
);

defparam ram16sdp_inst_320.INIT_0 = 16'h0000;
defparam ram16sdp_inst_320.INIT_1 = 16'h0000;
defparam ram16sdp_inst_320.INIT_2 = 16'h0000;
defparam ram16sdp_inst_320.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_321 (
    .DO(ram16sdp_inst_321_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_122),
    .CLK(clk)
);

defparam ram16sdp_inst_321.INIT_0 = 16'h0000;
defparam ram16sdp_inst_321.INIT_1 = 16'h0000;
defparam ram16sdp_inst_321.INIT_2 = 16'h0000;
defparam ram16sdp_inst_321.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_322 (
    .DO(ram16sdp_inst_322_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_122),
    .CLK(clk)
);

defparam ram16sdp_inst_322.INIT_0 = 16'h0000;
defparam ram16sdp_inst_322.INIT_1 = 16'h0000;
defparam ram16sdp_inst_322.INIT_2 = 16'h0000;
defparam ram16sdp_inst_322.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_323 (
    .DO(ram16sdp_inst_323_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_122),
    .CLK(clk)
);

defparam ram16sdp_inst_323.INIT_0 = 16'h0000;
defparam ram16sdp_inst_323.INIT_1 = 16'h0000;
defparam ram16sdp_inst_323.INIT_2 = 16'h0000;
defparam ram16sdp_inst_323.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_324 (
    .DO(ram16sdp_inst_324_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_122),
    .CLK(clk)
);

defparam ram16sdp_inst_324.INIT_0 = 16'h0000;
defparam ram16sdp_inst_324.INIT_1 = 16'h0000;
defparam ram16sdp_inst_324.INIT_2 = 16'h0000;
defparam ram16sdp_inst_324.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_325 (
    .DO(ram16sdp_inst_325_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_122),
    .CLK(clk)
);

defparam ram16sdp_inst_325.INIT_0 = 16'h0000;
defparam ram16sdp_inst_325.INIT_1 = 16'h0000;
defparam ram16sdp_inst_325.INIT_2 = 16'h0000;
defparam ram16sdp_inst_325.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_326 (
    .DO(ram16sdp_inst_326_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_122),
    .CLK(clk)
);

defparam ram16sdp_inst_326.INIT_0 = 16'h0000;
defparam ram16sdp_inst_326.INIT_1 = 16'h0000;
defparam ram16sdp_inst_326.INIT_2 = 16'h0000;
defparam ram16sdp_inst_326.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_327 (
    .DO(ram16sdp_inst_327_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_122),
    .CLK(clk)
);

defparam ram16sdp_inst_327.INIT_0 = 16'h0000;
defparam ram16sdp_inst_327.INIT_1 = 16'h0000;
defparam ram16sdp_inst_327.INIT_2 = 16'h0000;
defparam ram16sdp_inst_327.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_328 (
    .DO(ram16sdp_inst_328_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_125),
    .CLK(clk)
);

defparam ram16sdp_inst_328.INIT_0 = 16'h0000;
defparam ram16sdp_inst_328.INIT_1 = 16'h0000;
defparam ram16sdp_inst_328.INIT_2 = 16'h0000;
defparam ram16sdp_inst_328.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_329 (
    .DO(ram16sdp_inst_329_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_125),
    .CLK(clk)
);

defparam ram16sdp_inst_329.INIT_0 = 16'h0000;
defparam ram16sdp_inst_329.INIT_1 = 16'h0000;
defparam ram16sdp_inst_329.INIT_2 = 16'h0000;
defparam ram16sdp_inst_329.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_330 (
    .DO(ram16sdp_inst_330_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_125),
    .CLK(clk)
);

defparam ram16sdp_inst_330.INIT_0 = 16'h0000;
defparam ram16sdp_inst_330.INIT_1 = 16'h0000;
defparam ram16sdp_inst_330.INIT_2 = 16'h0000;
defparam ram16sdp_inst_330.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_331 (
    .DO(ram16sdp_inst_331_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_125),
    .CLK(clk)
);

defparam ram16sdp_inst_331.INIT_0 = 16'h0000;
defparam ram16sdp_inst_331.INIT_1 = 16'h0000;
defparam ram16sdp_inst_331.INIT_2 = 16'h0000;
defparam ram16sdp_inst_331.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_332 (
    .DO(ram16sdp_inst_332_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_125),
    .CLK(clk)
);

defparam ram16sdp_inst_332.INIT_0 = 16'h0000;
defparam ram16sdp_inst_332.INIT_1 = 16'h0000;
defparam ram16sdp_inst_332.INIT_2 = 16'h0000;
defparam ram16sdp_inst_332.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_333 (
    .DO(ram16sdp_inst_333_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_125),
    .CLK(clk)
);

defparam ram16sdp_inst_333.INIT_0 = 16'h0000;
defparam ram16sdp_inst_333.INIT_1 = 16'h0000;
defparam ram16sdp_inst_333.INIT_2 = 16'h0000;
defparam ram16sdp_inst_333.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_334 (
    .DO(ram16sdp_inst_334_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_125),
    .CLK(clk)
);

defparam ram16sdp_inst_334.INIT_0 = 16'h0000;
defparam ram16sdp_inst_334.INIT_1 = 16'h0000;
defparam ram16sdp_inst_334.INIT_2 = 16'h0000;
defparam ram16sdp_inst_334.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_335 (
    .DO(ram16sdp_inst_335_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_125),
    .CLK(clk)
);

defparam ram16sdp_inst_335.INIT_0 = 16'h0000;
defparam ram16sdp_inst_335.INIT_1 = 16'h0000;
defparam ram16sdp_inst_335.INIT_2 = 16'h0000;
defparam ram16sdp_inst_335.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_336 (
    .DO(ram16sdp_inst_336_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_128),
    .CLK(clk)
);

defparam ram16sdp_inst_336.INIT_0 = 16'h0000;
defparam ram16sdp_inst_336.INIT_1 = 16'h0000;
defparam ram16sdp_inst_336.INIT_2 = 16'h0000;
defparam ram16sdp_inst_336.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_337 (
    .DO(ram16sdp_inst_337_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_128),
    .CLK(clk)
);

defparam ram16sdp_inst_337.INIT_0 = 16'h0000;
defparam ram16sdp_inst_337.INIT_1 = 16'h0000;
defparam ram16sdp_inst_337.INIT_2 = 16'h0000;
defparam ram16sdp_inst_337.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_338 (
    .DO(ram16sdp_inst_338_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_128),
    .CLK(clk)
);

defparam ram16sdp_inst_338.INIT_0 = 16'h0000;
defparam ram16sdp_inst_338.INIT_1 = 16'h0000;
defparam ram16sdp_inst_338.INIT_2 = 16'h0000;
defparam ram16sdp_inst_338.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_339 (
    .DO(ram16sdp_inst_339_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_128),
    .CLK(clk)
);

defparam ram16sdp_inst_339.INIT_0 = 16'h0000;
defparam ram16sdp_inst_339.INIT_1 = 16'h0000;
defparam ram16sdp_inst_339.INIT_2 = 16'h0000;
defparam ram16sdp_inst_339.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_340 (
    .DO(ram16sdp_inst_340_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_128),
    .CLK(clk)
);

defparam ram16sdp_inst_340.INIT_0 = 16'h0000;
defparam ram16sdp_inst_340.INIT_1 = 16'h0000;
defparam ram16sdp_inst_340.INIT_2 = 16'h0000;
defparam ram16sdp_inst_340.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_341 (
    .DO(ram16sdp_inst_341_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_128),
    .CLK(clk)
);

defparam ram16sdp_inst_341.INIT_0 = 16'h0000;
defparam ram16sdp_inst_341.INIT_1 = 16'h0000;
defparam ram16sdp_inst_341.INIT_2 = 16'h0000;
defparam ram16sdp_inst_341.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_342 (
    .DO(ram16sdp_inst_342_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_128),
    .CLK(clk)
);

defparam ram16sdp_inst_342.INIT_0 = 16'h0000;
defparam ram16sdp_inst_342.INIT_1 = 16'h0000;
defparam ram16sdp_inst_342.INIT_2 = 16'h0000;
defparam ram16sdp_inst_342.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_343 (
    .DO(ram16sdp_inst_343_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_128),
    .CLK(clk)
);

defparam ram16sdp_inst_343.INIT_0 = 16'h0000;
defparam ram16sdp_inst_343.INIT_1 = 16'h0000;
defparam ram16sdp_inst_343.INIT_2 = 16'h0000;
defparam ram16sdp_inst_343.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_344 (
    .DO(ram16sdp_inst_344_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16sdp_inst_344.INIT_0 = 16'h0000;
defparam ram16sdp_inst_344.INIT_1 = 16'h0000;
defparam ram16sdp_inst_344.INIT_2 = 16'h0000;
defparam ram16sdp_inst_344.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_345 (
    .DO(ram16sdp_inst_345_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16sdp_inst_345.INIT_0 = 16'h0000;
defparam ram16sdp_inst_345.INIT_1 = 16'h0000;
defparam ram16sdp_inst_345.INIT_2 = 16'h0000;
defparam ram16sdp_inst_345.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_346 (
    .DO(ram16sdp_inst_346_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16sdp_inst_346.INIT_0 = 16'h0000;
defparam ram16sdp_inst_346.INIT_1 = 16'h0000;
defparam ram16sdp_inst_346.INIT_2 = 16'h0000;
defparam ram16sdp_inst_346.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_347 (
    .DO(ram16sdp_inst_347_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16sdp_inst_347.INIT_0 = 16'h0000;
defparam ram16sdp_inst_347.INIT_1 = 16'h0000;
defparam ram16sdp_inst_347.INIT_2 = 16'h0000;
defparam ram16sdp_inst_347.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_348 (
    .DO(ram16sdp_inst_348_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16sdp_inst_348.INIT_0 = 16'h0000;
defparam ram16sdp_inst_348.INIT_1 = 16'h0000;
defparam ram16sdp_inst_348.INIT_2 = 16'h0000;
defparam ram16sdp_inst_348.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_349 (
    .DO(ram16sdp_inst_349_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16sdp_inst_349.INIT_0 = 16'h0000;
defparam ram16sdp_inst_349.INIT_1 = 16'h0000;
defparam ram16sdp_inst_349.INIT_2 = 16'h0000;
defparam ram16sdp_inst_349.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_350 (
    .DO(ram16sdp_inst_350_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16sdp_inst_350.INIT_0 = 16'h0000;
defparam ram16sdp_inst_350.INIT_1 = 16'h0000;
defparam ram16sdp_inst_350.INIT_2 = 16'h0000;
defparam ram16sdp_inst_350.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_351 (
    .DO(ram16sdp_inst_351_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16sdp_inst_351.INIT_0 = 16'h0000;
defparam ram16sdp_inst_351.INIT_1 = 16'h0000;
defparam ram16sdp_inst_351.INIT_2 = 16'h0000;
defparam ram16sdp_inst_351.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_352 (
    .DO(ram16sdp_inst_352_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_134),
    .CLK(clk)
);

defparam ram16sdp_inst_352.INIT_0 = 16'h0000;
defparam ram16sdp_inst_352.INIT_1 = 16'h0000;
defparam ram16sdp_inst_352.INIT_2 = 16'h0000;
defparam ram16sdp_inst_352.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_353 (
    .DO(ram16sdp_inst_353_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_134),
    .CLK(clk)
);

defparam ram16sdp_inst_353.INIT_0 = 16'h0000;
defparam ram16sdp_inst_353.INIT_1 = 16'h0000;
defparam ram16sdp_inst_353.INIT_2 = 16'h0000;
defparam ram16sdp_inst_353.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_354 (
    .DO(ram16sdp_inst_354_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_134),
    .CLK(clk)
);

defparam ram16sdp_inst_354.INIT_0 = 16'h0000;
defparam ram16sdp_inst_354.INIT_1 = 16'h0000;
defparam ram16sdp_inst_354.INIT_2 = 16'h0000;
defparam ram16sdp_inst_354.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_355 (
    .DO(ram16sdp_inst_355_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_134),
    .CLK(clk)
);

defparam ram16sdp_inst_355.INIT_0 = 16'h0000;
defparam ram16sdp_inst_355.INIT_1 = 16'h0000;
defparam ram16sdp_inst_355.INIT_2 = 16'h0000;
defparam ram16sdp_inst_355.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_356 (
    .DO(ram16sdp_inst_356_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_134),
    .CLK(clk)
);

defparam ram16sdp_inst_356.INIT_0 = 16'h0000;
defparam ram16sdp_inst_356.INIT_1 = 16'h0000;
defparam ram16sdp_inst_356.INIT_2 = 16'h0000;
defparam ram16sdp_inst_356.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_357 (
    .DO(ram16sdp_inst_357_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_134),
    .CLK(clk)
);

defparam ram16sdp_inst_357.INIT_0 = 16'h0000;
defparam ram16sdp_inst_357.INIT_1 = 16'h0000;
defparam ram16sdp_inst_357.INIT_2 = 16'h0000;
defparam ram16sdp_inst_357.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_358 (
    .DO(ram16sdp_inst_358_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_134),
    .CLK(clk)
);

defparam ram16sdp_inst_358.INIT_0 = 16'h0000;
defparam ram16sdp_inst_358.INIT_1 = 16'h0000;
defparam ram16sdp_inst_358.INIT_2 = 16'h0000;
defparam ram16sdp_inst_358.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_359 (
    .DO(ram16sdp_inst_359_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_134),
    .CLK(clk)
);

defparam ram16sdp_inst_359.INIT_0 = 16'h0000;
defparam ram16sdp_inst_359.INIT_1 = 16'h0000;
defparam ram16sdp_inst_359.INIT_2 = 16'h0000;
defparam ram16sdp_inst_359.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_360 (
    .DO(ram16sdp_inst_360_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_137),
    .CLK(clk)
);

defparam ram16sdp_inst_360.INIT_0 = 16'h0000;
defparam ram16sdp_inst_360.INIT_1 = 16'h0000;
defparam ram16sdp_inst_360.INIT_2 = 16'h0000;
defparam ram16sdp_inst_360.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_361 (
    .DO(ram16sdp_inst_361_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_137),
    .CLK(clk)
);

defparam ram16sdp_inst_361.INIT_0 = 16'h0000;
defparam ram16sdp_inst_361.INIT_1 = 16'h0000;
defparam ram16sdp_inst_361.INIT_2 = 16'h0000;
defparam ram16sdp_inst_361.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_362 (
    .DO(ram16sdp_inst_362_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_137),
    .CLK(clk)
);

defparam ram16sdp_inst_362.INIT_0 = 16'h0000;
defparam ram16sdp_inst_362.INIT_1 = 16'h0000;
defparam ram16sdp_inst_362.INIT_2 = 16'h0000;
defparam ram16sdp_inst_362.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_363 (
    .DO(ram16sdp_inst_363_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_137),
    .CLK(clk)
);

defparam ram16sdp_inst_363.INIT_0 = 16'h0000;
defparam ram16sdp_inst_363.INIT_1 = 16'h0000;
defparam ram16sdp_inst_363.INIT_2 = 16'h0000;
defparam ram16sdp_inst_363.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_364 (
    .DO(ram16sdp_inst_364_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_137),
    .CLK(clk)
);

defparam ram16sdp_inst_364.INIT_0 = 16'h0000;
defparam ram16sdp_inst_364.INIT_1 = 16'h0000;
defparam ram16sdp_inst_364.INIT_2 = 16'h0000;
defparam ram16sdp_inst_364.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_365 (
    .DO(ram16sdp_inst_365_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_137),
    .CLK(clk)
);

defparam ram16sdp_inst_365.INIT_0 = 16'h0000;
defparam ram16sdp_inst_365.INIT_1 = 16'h0000;
defparam ram16sdp_inst_365.INIT_2 = 16'h0000;
defparam ram16sdp_inst_365.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_366 (
    .DO(ram16sdp_inst_366_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_137),
    .CLK(clk)
);

defparam ram16sdp_inst_366.INIT_0 = 16'h0000;
defparam ram16sdp_inst_366.INIT_1 = 16'h0000;
defparam ram16sdp_inst_366.INIT_2 = 16'h0000;
defparam ram16sdp_inst_366.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_367 (
    .DO(ram16sdp_inst_367_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_137),
    .CLK(clk)
);

defparam ram16sdp_inst_367.INIT_0 = 16'h0000;
defparam ram16sdp_inst_367.INIT_1 = 16'h0000;
defparam ram16sdp_inst_367.INIT_2 = 16'h0000;
defparam ram16sdp_inst_367.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_368 (
    .DO(ram16sdp_inst_368_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_140),
    .CLK(clk)
);

defparam ram16sdp_inst_368.INIT_0 = 16'h0000;
defparam ram16sdp_inst_368.INIT_1 = 16'h0000;
defparam ram16sdp_inst_368.INIT_2 = 16'h0000;
defparam ram16sdp_inst_368.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_369 (
    .DO(ram16sdp_inst_369_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_140),
    .CLK(clk)
);

defparam ram16sdp_inst_369.INIT_0 = 16'h0000;
defparam ram16sdp_inst_369.INIT_1 = 16'h0000;
defparam ram16sdp_inst_369.INIT_2 = 16'h0000;
defparam ram16sdp_inst_369.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_370 (
    .DO(ram16sdp_inst_370_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_140),
    .CLK(clk)
);

defparam ram16sdp_inst_370.INIT_0 = 16'h0000;
defparam ram16sdp_inst_370.INIT_1 = 16'h0000;
defparam ram16sdp_inst_370.INIT_2 = 16'h0000;
defparam ram16sdp_inst_370.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_371 (
    .DO(ram16sdp_inst_371_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_140),
    .CLK(clk)
);

defparam ram16sdp_inst_371.INIT_0 = 16'h0000;
defparam ram16sdp_inst_371.INIT_1 = 16'h0000;
defparam ram16sdp_inst_371.INIT_2 = 16'h0000;
defparam ram16sdp_inst_371.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_372 (
    .DO(ram16sdp_inst_372_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_140),
    .CLK(clk)
);

defparam ram16sdp_inst_372.INIT_0 = 16'h0000;
defparam ram16sdp_inst_372.INIT_1 = 16'h0000;
defparam ram16sdp_inst_372.INIT_2 = 16'h0000;
defparam ram16sdp_inst_372.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_373 (
    .DO(ram16sdp_inst_373_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_140),
    .CLK(clk)
);

defparam ram16sdp_inst_373.INIT_0 = 16'h0000;
defparam ram16sdp_inst_373.INIT_1 = 16'h0000;
defparam ram16sdp_inst_373.INIT_2 = 16'h0000;
defparam ram16sdp_inst_373.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_374 (
    .DO(ram16sdp_inst_374_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_140),
    .CLK(clk)
);

defparam ram16sdp_inst_374.INIT_0 = 16'h0000;
defparam ram16sdp_inst_374.INIT_1 = 16'h0000;
defparam ram16sdp_inst_374.INIT_2 = 16'h0000;
defparam ram16sdp_inst_374.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_375 (
    .DO(ram16sdp_inst_375_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_140),
    .CLK(clk)
);

defparam ram16sdp_inst_375.INIT_0 = 16'h0000;
defparam ram16sdp_inst_375.INIT_1 = 16'h0000;
defparam ram16sdp_inst_375.INIT_2 = 16'h0000;
defparam ram16sdp_inst_375.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_376 (
    .DO(ram16sdp_inst_376_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16sdp_inst_376.INIT_0 = 16'h0000;
defparam ram16sdp_inst_376.INIT_1 = 16'h0000;
defparam ram16sdp_inst_376.INIT_2 = 16'h0000;
defparam ram16sdp_inst_376.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_377 (
    .DO(ram16sdp_inst_377_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16sdp_inst_377.INIT_0 = 16'h0000;
defparam ram16sdp_inst_377.INIT_1 = 16'h0000;
defparam ram16sdp_inst_377.INIT_2 = 16'h0000;
defparam ram16sdp_inst_377.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_378 (
    .DO(ram16sdp_inst_378_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16sdp_inst_378.INIT_0 = 16'h0000;
defparam ram16sdp_inst_378.INIT_1 = 16'h0000;
defparam ram16sdp_inst_378.INIT_2 = 16'h0000;
defparam ram16sdp_inst_378.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_379 (
    .DO(ram16sdp_inst_379_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16sdp_inst_379.INIT_0 = 16'h0000;
defparam ram16sdp_inst_379.INIT_1 = 16'h0000;
defparam ram16sdp_inst_379.INIT_2 = 16'h0000;
defparam ram16sdp_inst_379.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_380 (
    .DO(ram16sdp_inst_380_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16sdp_inst_380.INIT_0 = 16'h0000;
defparam ram16sdp_inst_380.INIT_1 = 16'h0000;
defparam ram16sdp_inst_380.INIT_2 = 16'h0000;
defparam ram16sdp_inst_380.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_381 (
    .DO(ram16sdp_inst_381_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16sdp_inst_381.INIT_0 = 16'h0000;
defparam ram16sdp_inst_381.INIT_1 = 16'h0000;
defparam ram16sdp_inst_381.INIT_2 = 16'h0000;
defparam ram16sdp_inst_381.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_382 (
    .DO(ram16sdp_inst_382_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16sdp_inst_382.INIT_0 = 16'h0000;
defparam ram16sdp_inst_382.INIT_1 = 16'h0000;
defparam ram16sdp_inst_382.INIT_2 = 16'h0000;
defparam ram16sdp_inst_382.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_383 (
    .DO(ram16sdp_inst_383_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16sdp_inst_383.INIT_0 = 16'h0000;
defparam ram16sdp_inst_383.INIT_1 = 16'h0000;
defparam ram16sdp_inst_383.INIT_2 = 16'h0000;
defparam ram16sdp_inst_383.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_384 (
    .DO(ram16sdp_inst_384_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_146),
    .CLK(clk)
);

defparam ram16sdp_inst_384.INIT_0 = 16'h0000;
defparam ram16sdp_inst_384.INIT_1 = 16'h0000;
defparam ram16sdp_inst_384.INIT_2 = 16'h0000;
defparam ram16sdp_inst_384.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_385 (
    .DO(ram16sdp_inst_385_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_146),
    .CLK(clk)
);

defparam ram16sdp_inst_385.INIT_0 = 16'h0000;
defparam ram16sdp_inst_385.INIT_1 = 16'h0000;
defparam ram16sdp_inst_385.INIT_2 = 16'h0000;
defparam ram16sdp_inst_385.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_386 (
    .DO(ram16sdp_inst_386_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_146),
    .CLK(clk)
);

defparam ram16sdp_inst_386.INIT_0 = 16'h0000;
defparam ram16sdp_inst_386.INIT_1 = 16'h0000;
defparam ram16sdp_inst_386.INIT_2 = 16'h0000;
defparam ram16sdp_inst_386.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_387 (
    .DO(ram16sdp_inst_387_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_146),
    .CLK(clk)
);

defparam ram16sdp_inst_387.INIT_0 = 16'h0000;
defparam ram16sdp_inst_387.INIT_1 = 16'h0000;
defparam ram16sdp_inst_387.INIT_2 = 16'h0000;
defparam ram16sdp_inst_387.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_388 (
    .DO(ram16sdp_inst_388_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_146),
    .CLK(clk)
);

defparam ram16sdp_inst_388.INIT_0 = 16'h0000;
defparam ram16sdp_inst_388.INIT_1 = 16'h0000;
defparam ram16sdp_inst_388.INIT_2 = 16'h0000;
defparam ram16sdp_inst_388.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_389 (
    .DO(ram16sdp_inst_389_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_146),
    .CLK(clk)
);

defparam ram16sdp_inst_389.INIT_0 = 16'h0000;
defparam ram16sdp_inst_389.INIT_1 = 16'h0000;
defparam ram16sdp_inst_389.INIT_2 = 16'h0000;
defparam ram16sdp_inst_389.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_390 (
    .DO(ram16sdp_inst_390_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_146),
    .CLK(clk)
);

defparam ram16sdp_inst_390.INIT_0 = 16'h0000;
defparam ram16sdp_inst_390.INIT_1 = 16'h0000;
defparam ram16sdp_inst_390.INIT_2 = 16'h0000;
defparam ram16sdp_inst_390.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_391 (
    .DO(ram16sdp_inst_391_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_146),
    .CLK(clk)
);

defparam ram16sdp_inst_391.INIT_0 = 16'h0000;
defparam ram16sdp_inst_391.INIT_1 = 16'h0000;
defparam ram16sdp_inst_391.INIT_2 = 16'h0000;
defparam ram16sdp_inst_391.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_392 (
    .DO(ram16sdp_inst_392_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_149),
    .CLK(clk)
);

defparam ram16sdp_inst_392.INIT_0 = 16'h0000;
defparam ram16sdp_inst_392.INIT_1 = 16'h0000;
defparam ram16sdp_inst_392.INIT_2 = 16'h0000;
defparam ram16sdp_inst_392.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_393 (
    .DO(ram16sdp_inst_393_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_149),
    .CLK(clk)
);

defparam ram16sdp_inst_393.INIT_0 = 16'h0000;
defparam ram16sdp_inst_393.INIT_1 = 16'h0000;
defparam ram16sdp_inst_393.INIT_2 = 16'h0000;
defparam ram16sdp_inst_393.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_394 (
    .DO(ram16sdp_inst_394_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_149),
    .CLK(clk)
);

defparam ram16sdp_inst_394.INIT_0 = 16'h0000;
defparam ram16sdp_inst_394.INIT_1 = 16'h0000;
defparam ram16sdp_inst_394.INIT_2 = 16'h0000;
defparam ram16sdp_inst_394.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_395 (
    .DO(ram16sdp_inst_395_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_149),
    .CLK(clk)
);

defparam ram16sdp_inst_395.INIT_0 = 16'h0000;
defparam ram16sdp_inst_395.INIT_1 = 16'h0000;
defparam ram16sdp_inst_395.INIT_2 = 16'h0000;
defparam ram16sdp_inst_395.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_396 (
    .DO(ram16sdp_inst_396_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_149),
    .CLK(clk)
);

defparam ram16sdp_inst_396.INIT_0 = 16'h0000;
defparam ram16sdp_inst_396.INIT_1 = 16'h0000;
defparam ram16sdp_inst_396.INIT_2 = 16'h0000;
defparam ram16sdp_inst_396.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_397 (
    .DO(ram16sdp_inst_397_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_149),
    .CLK(clk)
);

defparam ram16sdp_inst_397.INIT_0 = 16'h0000;
defparam ram16sdp_inst_397.INIT_1 = 16'h0000;
defparam ram16sdp_inst_397.INIT_2 = 16'h0000;
defparam ram16sdp_inst_397.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_398 (
    .DO(ram16sdp_inst_398_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_149),
    .CLK(clk)
);

defparam ram16sdp_inst_398.INIT_0 = 16'h0000;
defparam ram16sdp_inst_398.INIT_1 = 16'h0000;
defparam ram16sdp_inst_398.INIT_2 = 16'h0000;
defparam ram16sdp_inst_398.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_399 (
    .DO(ram16sdp_inst_399_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_149),
    .CLK(clk)
);

defparam ram16sdp_inst_399.INIT_0 = 16'h0000;
defparam ram16sdp_inst_399.INIT_1 = 16'h0000;
defparam ram16sdp_inst_399.INIT_2 = 16'h0000;
defparam ram16sdp_inst_399.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_400 (
    .DO(ram16sdp_inst_400_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_152),
    .CLK(clk)
);

defparam ram16sdp_inst_400.INIT_0 = 16'h0000;
defparam ram16sdp_inst_400.INIT_1 = 16'h0000;
defparam ram16sdp_inst_400.INIT_2 = 16'h0000;
defparam ram16sdp_inst_400.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_401 (
    .DO(ram16sdp_inst_401_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_152),
    .CLK(clk)
);

defparam ram16sdp_inst_401.INIT_0 = 16'h0000;
defparam ram16sdp_inst_401.INIT_1 = 16'h0000;
defparam ram16sdp_inst_401.INIT_2 = 16'h0000;
defparam ram16sdp_inst_401.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_402 (
    .DO(ram16sdp_inst_402_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_152),
    .CLK(clk)
);

defparam ram16sdp_inst_402.INIT_0 = 16'h0000;
defparam ram16sdp_inst_402.INIT_1 = 16'h0000;
defparam ram16sdp_inst_402.INIT_2 = 16'h0000;
defparam ram16sdp_inst_402.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_403 (
    .DO(ram16sdp_inst_403_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_152),
    .CLK(clk)
);

defparam ram16sdp_inst_403.INIT_0 = 16'h0000;
defparam ram16sdp_inst_403.INIT_1 = 16'h0000;
defparam ram16sdp_inst_403.INIT_2 = 16'h0000;
defparam ram16sdp_inst_403.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_404 (
    .DO(ram16sdp_inst_404_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_152),
    .CLK(clk)
);

defparam ram16sdp_inst_404.INIT_0 = 16'h0000;
defparam ram16sdp_inst_404.INIT_1 = 16'h0000;
defparam ram16sdp_inst_404.INIT_2 = 16'h0000;
defparam ram16sdp_inst_404.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_405 (
    .DO(ram16sdp_inst_405_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_152),
    .CLK(clk)
);

defparam ram16sdp_inst_405.INIT_0 = 16'h0000;
defparam ram16sdp_inst_405.INIT_1 = 16'h0000;
defparam ram16sdp_inst_405.INIT_2 = 16'h0000;
defparam ram16sdp_inst_405.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_406 (
    .DO(ram16sdp_inst_406_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_152),
    .CLK(clk)
);

defparam ram16sdp_inst_406.INIT_0 = 16'h0000;
defparam ram16sdp_inst_406.INIT_1 = 16'h0000;
defparam ram16sdp_inst_406.INIT_2 = 16'h0000;
defparam ram16sdp_inst_406.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_407 (
    .DO(ram16sdp_inst_407_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_152),
    .CLK(clk)
);

defparam ram16sdp_inst_407.INIT_0 = 16'h0000;
defparam ram16sdp_inst_407.INIT_1 = 16'h0000;
defparam ram16sdp_inst_407.INIT_2 = 16'h0000;
defparam ram16sdp_inst_407.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_408 (
    .DO(ram16sdp_inst_408_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16sdp_inst_408.INIT_0 = 16'h0000;
defparam ram16sdp_inst_408.INIT_1 = 16'h0000;
defparam ram16sdp_inst_408.INIT_2 = 16'h0000;
defparam ram16sdp_inst_408.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_409 (
    .DO(ram16sdp_inst_409_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16sdp_inst_409.INIT_0 = 16'h0000;
defparam ram16sdp_inst_409.INIT_1 = 16'h0000;
defparam ram16sdp_inst_409.INIT_2 = 16'h0000;
defparam ram16sdp_inst_409.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_410 (
    .DO(ram16sdp_inst_410_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16sdp_inst_410.INIT_0 = 16'h0000;
defparam ram16sdp_inst_410.INIT_1 = 16'h0000;
defparam ram16sdp_inst_410.INIT_2 = 16'h0000;
defparam ram16sdp_inst_410.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_411 (
    .DO(ram16sdp_inst_411_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16sdp_inst_411.INIT_0 = 16'h0000;
defparam ram16sdp_inst_411.INIT_1 = 16'h0000;
defparam ram16sdp_inst_411.INIT_2 = 16'h0000;
defparam ram16sdp_inst_411.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_412 (
    .DO(ram16sdp_inst_412_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16sdp_inst_412.INIT_0 = 16'h0000;
defparam ram16sdp_inst_412.INIT_1 = 16'h0000;
defparam ram16sdp_inst_412.INIT_2 = 16'h0000;
defparam ram16sdp_inst_412.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_413 (
    .DO(ram16sdp_inst_413_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16sdp_inst_413.INIT_0 = 16'h0000;
defparam ram16sdp_inst_413.INIT_1 = 16'h0000;
defparam ram16sdp_inst_413.INIT_2 = 16'h0000;
defparam ram16sdp_inst_413.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_414 (
    .DO(ram16sdp_inst_414_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16sdp_inst_414.INIT_0 = 16'h0000;
defparam ram16sdp_inst_414.INIT_1 = 16'h0000;
defparam ram16sdp_inst_414.INIT_2 = 16'h0000;
defparam ram16sdp_inst_414.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_415 (
    .DO(ram16sdp_inst_415_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16sdp_inst_415.INIT_0 = 16'h0000;
defparam ram16sdp_inst_415.INIT_1 = 16'h0000;
defparam ram16sdp_inst_415.INIT_2 = 16'h0000;
defparam ram16sdp_inst_415.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_416 (
    .DO(ram16sdp_inst_416_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_158),
    .CLK(clk)
);

defparam ram16sdp_inst_416.INIT_0 = 16'h0000;
defparam ram16sdp_inst_416.INIT_1 = 16'h0000;
defparam ram16sdp_inst_416.INIT_2 = 16'h0000;
defparam ram16sdp_inst_416.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_417 (
    .DO(ram16sdp_inst_417_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_158),
    .CLK(clk)
);

defparam ram16sdp_inst_417.INIT_0 = 16'h0000;
defparam ram16sdp_inst_417.INIT_1 = 16'h0000;
defparam ram16sdp_inst_417.INIT_2 = 16'h0000;
defparam ram16sdp_inst_417.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_418 (
    .DO(ram16sdp_inst_418_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_158),
    .CLK(clk)
);

defparam ram16sdp_inst_418.INIT_0 = 16'h0000;
defparam ram16sdp_inst_418.INIT_1 = 16'h0000;
defparam ram16sdp_inst_418.INIT_2 = 16'h0000;
defparam ram16sdp_inst_418.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_419 (
    .DO(ram16sdp_inst_419_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_158),
    .CLK(clk)
);

defparam ram16sdp_inst_419.INIT_0 = 16'h0000;
defparam ram16sdp_inst_419.INIT_1 = 16'h0000;
defparam ram16sdp_inst_419.INIT_2 = 16'h0000;
defparam ram16sdp_inst_419.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_420 (
    .DO(ram16sdp_inst_420_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_158),
    .CLK(clk)
);

defparam ram16sdp_inst_420.INIT_0 = 16'h0000;
defparam ram16sdp_inst_420.INIT_1 = 16'h0000;
defparam ram16sdp_inst_420.INIT_2 = 16'h0000;
defparam ram16sdp_inst_420.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_421 (
    .DO(ram16sdp_inst_421_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_158),
    .CLK(clk)
);

defparam ram16sdp_inst_421.INIT_0 = 16'h0000;
defparam ram16sdp_inst_421.INIT_1 = 16'h0000;
defparam ram16sdp_inst_421.INIT_2 = 16'h0000;
defparam ram16sdp_inst_421.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_422 (
    .DO(ram16sdp_inst_422_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_158),
    .CLK(clk)
);

defparam ram16sdp_inst_422.INIT_0 = 16'h0000;
defparam ram16sdp_inst_422.INIT_1 = 16'h0000;
defparam ram16sdp_inst_422.INIT_2 = 16'h0000;
defparam ram16sdp_inst_422.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_423 (
    .DO(ram16sdp_inst_423_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_158),
    .CLK(clk)
);

defparam ram16sdp_inst_423.INIT_0 = 16'h0000;
defparam ram16sdp_inst_423.INIT_1 = 16'h0000;
defparam ram16sdp_inst_423.INIT_2 = 16'h0000;
defparam ram16sdp_inst_423.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_424 (
    .DO(ram16sdp_inst_424_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_161),
    .CLK(clk)
);

defparam ram16sdp_inst_424.INIT_0 = 16'h0000;
defparam ram16sdp_inst_424.INIT_1 = 16'h0000;
defparam ram16sdp_inst_424.INIT_2 = 16'h0000;
defparam ram16sdp_inst_424.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_425 (
    .DO(ram16sdp_inst_425_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_161),
    .CLK(clk)
);

defparam ram16sdp_inst_425.INIT_0 = 16'h0000;
defparam ram16sdp_inst_425.INIT_1 = 16'h0000;
defparam ram16sdp_inst_425.INIT_2 = 16'h0000;
defparam ram16sdp_inst_425.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_426 (
    .DO(ram16sdp_inst_426_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_161),
    .CLK(clk)
);

defparam ram16sdp_inst_426.INIT_0 = 16'h0000;
defparam ram16sdp_inst_426.INIT_1 = 16'h0000;
defparam ram16sdp_inst_426.INIT_2 = 16'h0000;
defparam ram16sdp_inst_426.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_427 (
    .DO(ram16sdp_inst_427_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_161),
    .CLK(clk)
);

defparam ram16sdp_inst_427.INIT_0 = 16'h0000;
defparam ram16sdp_inst_427.INIT_1 = 16'h0000;
defparam ram16sdp_inst_427.INIT_2 = 16'h0000;
defparam ram16sdp_inst_427.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_428 (
    .DO(ram16sdp_inst_428_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_161),
    .CLK(clk)
);

defparam ram16sdp_inst_428.INIT_0 = 16'h0000;
defparam ram16sdp_inst_428.INIT_1 = 16'h0000;
defparam ram16sdp_inst_428.INIT_2 = 16'h0000;
defparam ram16sdp_inst_428.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_429 (
    .DO(ram16sdp_inst_429_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_161),
    .CLK(clk)
);

defparam ram16sdp_inst_429.INIT_0 = 16'h0000;
defparam ram16sdp_inst_429.INIT_1 = 16'h0000;
defparam ram16sdp_inst_429.INIT_2 = 16'h0000;
defparam ram16sdp_inst_429.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_430 (
    .DO(ram16sdp_inst_430_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_161),
    .CLK(clk)
);

defparam ram16sdp_inst_430.INIT_0 = 16'h0000;
defparam ram16sdp_inst_430.INIT_1 = 16'h0000;
defparam ram16sdp_inst_430.INIT_2 = 16'h0000;
defparam ram16sdp_inst_430.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_431 (
    .DO(ram16sdp_inst_431_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_161),
    .CLK(clk)
);

defparam ram16sdp_inst_431.INIT_0 = 16'h0000;
defparam ram16sdp_inst_431.INIT_1 = 16'h0000;
defparam ram16sdp_inst_431.INIT_2 = 16'h0000;
defparam ram16sdp_inst_431.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_432 (
    .DO(ram16sdp_inst_432_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_164),
    .CLK(clk)
);

defparam ram16sdp_inst_432.INIT_0 = 16'h0000;
defparam ram16sdp_inst_432.INIT_1 = 16'h0000;
defparam ram16sdp_inst_432.INIT_2 = 16'h0000;
defparam ram16sdp_inst_432.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_433 (
    .DO(ram16sdp_inst_433_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_164),
    .CLK(clk)
);

defparam ram16sdp_inst_433.INIT_0 = 16'h0000;
defparam ram16sdp_inst_433.INIT_1 = 16'h0000;
defparam ram16sdp_inst_433.INIT_2 = 16'h0000;
defparam ram16sdp_inst_433.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_434 (
    .DO(ram16sdp_inst_434_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_164),
    .CLK(clk)
);

defparam ram16sdp_inst_434.INIT_0 = 16'h0000;
defparam ram16sdp_inst_434.INIT_1 = 16'h0000;
defparam ram16sdp_inst_434.INIT_2 = 16'h0000;
defparam ram16sdp_inst_434.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_435 (
    .DO(ram16sdp_inst_435_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_164),
    .CLK(clk)
);

defparam ram16sdp_inst_435.INIT_0 = 16'h0000;
defparam ram16sdp_inst_435.INIT_1 = 16'h0000;
defparam ram16sdp_inst_435.INIT_2 = 16'h0000;
defparam ram16sdp_inst_435.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_436 (
    .DO(ram16sdp_inst_436_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_164),
    .CLK(clk)
);

defparam ram16sdp_inst_436.INIT_0 = 16'h0000;
defparam ram16sdp_inst_436.INIT_1 = 16'h0000;
defparam ram16sdp_inst_436.INIT_2 = 16'h0000;
defparam ram16sdp_inst_436.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_437 (
    .DO(ram16sdp_inst_437_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_164),
    .CLK(clk)
);

defparam ram16sdp_inst_437.INIT_0 = 16'h0000;
defparam ram16sdp_inst_437.INIT_1 = 16'h0000;
defparam ram16sdp_inst_437.INIT_2 = 16'h0000;
defparam ram16sdp_inst_437.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_438 (
    .DO(ram16sdp_inst_438_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_164),
    .CLK(clk)
);

defparam ram16sdp_inst_438.INIT_0 = 16'h0000;
defparam ram16sdp_inst_438.INIT_1 = 16'h0000;
defparam ram16sdp_inst_438.INIT_2 = 16'h0000;
defparam ram16sdp_inst_438.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_439 (
    .DO(ram16sdp_inst_439_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_164),
    .CLK(clk)
);

defparam ram16sdp_inst_439.INIT_0 = 16'h0000;
defparam ram16sdp_inst_439.INIT_1 = 16'h0000;
defparam ram16sdp_inst_439.INIT_2 = 16'h0000;
defparam ram16sdp_inst_439.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_440 (
    .DO(ram16sdp_inst_440_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16sdp_inst_440.INIT_0 = 16'h0000;
defparam ram16sdp_inst_440.INIT_1 = 16'h0000;
defparam ram16sdp_inst_440.INIT_2 = 16'h0000;
defparam ram16sdp_inst_440.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_441 (
    .DO(ram16sdp_inst_441_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16sdp_inst_441.INIT_0 = 16'h0000;
defparam ram16sdp_inst_441.INIT_1 = 16'h0000;
defparam ram16sdp_inst_441.INIT_2 = 16'h0000;
defparam ram16sdp_inst_441.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_442 (
    .DO(ram16sdp_inst_442_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16sdp_inst_442.INIT_0 = 16'h0000;
defparam ram16sdp_inst_442.INIT_1 = 16'h0000;
defparam ram16sdp_inst_442.INIT_2 = 16'h0000;
defparam ram16sdp_inst_442.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_443 (
    .DO(ram16sdp_inst_443_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16sdp_inst_443.INIT_0 = 16'h0000;
defparam ram16sdp_inst_443.INIT_1 = 16'h0000;
defparam ram16sdp_inst_443.INIT_2 = 16'h0000;
defparam ram16sdp_inst_443.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_444 (
    .DO(ram16sdp_inst_444_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16sdp_inst_444.INIT_0 = 16'h0000;
defparam ram16sdp_inst_444.INIT_1 = 16'h0000;
defparam ram16sdp_inst_444.INIT_2 = 16'h0000;
defparam ram16sdp_inst_444.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_445 (
    .DO(ram16sdp_inst_445_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16sdp_inst_445.INIT_0 = 16'h0000;
defparam ram16sdp_inst_445.INIT_1 = 16'h0000;
defparam ram16sdp_inst_445.INIT_2 = 16'h0000;
defparam ram16sdp_inst_445.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_446 (
    .DO(ram16sdp_inst_446_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16sdp_inst_446.INIT_0 = 16'h0000;
defparam ram16sdp_inst_446.INIT_1 = 16'h0000;
defparam ram16sdp_inst_446.INIT_2 = 16'h0000;
defparam ram16sdp_inst_446.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_447 (
    .DO(ram16sdp_inst_447_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16sdp_inst_447.INIT_0 = 16'h0000;
defparam ram16sdp_inst_447.INIT_1 = 16'h0000;
defparam ram16sdp_inst_447.INIT_2 = 16'h0000;
defparam ram16sdp_inst_447.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_448 (
    .DO(ram16sdp_inst_448_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_170),
    .CLK(clk)
);

defparam ram16sdp_inst_448.INIT_0 = 16'h0000;
defparam ram16sdp_inst_448.INIT_1 = 16'h0000;
defparam ram16sdp_inst_448.INIT_2 = 16'h0000;
defparam ram16sdp_inst_448.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_449 (
    .DO(ram16sdp_inst_449_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_170),
    .CLK(clk)
);

defparam ram16sdp_inst_449.INIT_0 = 16'h0000;
defparam ram16sdp_inst_449.INIT_1 = 16'h0000;
defparam ram16sdp_inst_449.INIT_2 = 16'h0000;
defparam ram16sdp_inst_449.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_450 (
    .DO(ram16sdp_inst_450_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_170),
    .CLK(clk)
);

defparam ram16sdp_inst_450.INIT_0 = 16'h0000;
defparam ram16sdp_inst_450.INIT_1 = 16'h0000;
defparam ram16sdp_inst_450.INIT_2 = 16'h0000;
defparam ram16sdp_inst_450.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_451 (
    .DO(ram16sdp_inst_451_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_170),
    .CLK(clk)
);

defparam ram16sdp_inst_451.INIT_0 = 16'h0000;
defparam ram16sdp_inst_451.INIT_1 = 16'h0000;
defparam ram16sdp_inst_451.INIT_2 = 16'h0000;
defparam ram16sdp_inst_451.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_452 (
    .DO(ram16sdp_inst_452_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_170),
    .CLK(clk)
);

defparam ram16sdp_inst_452.INIT_0 = 16'h0000;
defparam ram16sdp_inst_452.INIT_1 = 16'h0000;
defparam ram16sdp_inst_452.INIT_2 = 16'h0000;
defparam ram16sdp_inst_452.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_453 (
    .DO(ram16sdp_inst_453_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_170),
    .CLK(clk)
);

defparam ram16sdp_inst_453.INIT_0 = 16'h0000;
defparam ram16sdp_inst_453.INIT_1 = 16'h0000;
defparam ram16sdp_inst_453.INIT_2 = 16'h0000;
defparam ram16sdp_inst_453.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_454 (
    .DO(ram16sdp_inst_454_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_170),
    .CLK(clk)
);

defparam ram16sdp_inst_454.INIT_0 = 16'h0000;
defparam ram16sdp_inst_454.INIT_1 = 16'h0000;
defparam ram16sdp_inst_454.INIT_2 = 16'h0000;
defparam ram16sdp_inst_454.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_455 (
    .DO(ram16sdp_inst_455_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_170),
    .CLK(clk)
);

defparam ram16sdp_inst_455.INIT_0 = 16'h0000;
defparam ram16sdp_inst_455.INIT_1 = 16'h0000;
defparam ram16sdp_inst_455.INIT_2 = 16'h0000;
defparam ram16sdp_inst_455.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_456 (
    .DO(ram16sdp_inst_456_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_173),
    .CLK(clk)
);

defparam ram16sdp_inst_456.INIT_0 = 16'h0000;
defparam ram16sdp_inst_456.INIT_1 = 16'h0000;
defparam ram16sdp_inst_456.INIT_2 = 16'h0000;
defparam ram16sdp_inst_456.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_457 (
    .DO(ram16sdp_inst_457_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_173),
    .CLK(clk)
);

defparam ram16sdp_inst_457.INIT_0 = 16'h0000;
defparam ram16sdp_inst_457.INIT_1 = 16'h0000;
defparam ram16sdp_inst_457.INIT_2 = 16'h0000;
defparam ram16sdp_inst_457.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_458 (
    .DO(ram16sdp_inst_458_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_173),
    .CLK(clk)
);

defparam ram16sdp_inst_458.INIT_0 = 16'h0000;
defparam ram16sdp_inst_458.INIT_1 = 16'h0000;
defparam ram16sdp_inst_458.INIT_2 = 16'h0000;
defparam ram16sdp_inst_458.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_459 (
    .DO(ram16sdp_inst_459_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_173),
    .CLK(clk)
);

defparam ram16sdp_inst_459.INIT_0 = 16'h0000;
defparam ram16sdp_inst_459.INIT_1 = 16'h0000;
defparam ram16sdp_inst_459.INIT_2 = 16'h0000;
defparam ram16sdp_inst_459.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_460 (
    .DO(ram16sdp_inst_460_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_173),
    .CLK(clk)
);

defparam ram16sdp_inst_460.INIT_0 = 16'h0000;
defparam ram16sdp_inst_460.INIT_1 = 16'h0000;
defparam ram16sdp_inst_460.INIT_2 = 16'h0000;
defparam ram16sdp_inst_460.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_461 (
    .DO(ram16sdp_inst_461_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_173),
    .CLK(clk)
);

defparam ram16sdp_inst_461.INIT_0 = 16'h0000;
defparam ram16sdp_inst_461.INIT_1 = 16'h0000;
defparam ram16sdp_inst_461.INIT_2 = 16'h0000;
defparam ram16sdp_inst_461.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_462 (
    .DO(ram16sdp_inst_462_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_173),
    .CLK(clk)
);

defparam ram16sdp_inst_462.INIT_0 = 16'h0000;
defparam ram16sdp_inst_462.INIT_1 = 16'h0000;
defparam ram16sdp_inst_462.INIT_2 = 16'h0000;
defparam ram16sdp_inst_462.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_463 (
    .DO(ram16sdp_inst_463_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_173),
    .CLK(clk)
);

defparam ram16sdp_inst_463.INIT_0 = 16'h0000;
defparam ram16sdp_inst_463.INIT_1 = 16'h0000;
defparam ram16sdp_inst_463.INIT_2 = 16'h0000;
defparam ram16sdp_inst_463.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_464 (
    .DO(ram16sdp_inst_464_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_176),
    .CLK(clk)
);

defparam ram16sdp_inst_464.INIT_0 = 16'h0000;
defparam ram16sdp_inst_464.INIT_1 = 16'h0000;
defparam ram16sdp_inst_464.INIT_2 = 16'h0000;
defparam ram16sdp_inst_464.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_465 (
    .DO(ram16sdp_inst_465_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_176),
    .CLK(clk)
);

defparam ram16sdp_inst_465.INIT_0 = 16'h0000;
defparam ram16sdp_inst_465.INIT_1 = 16'h0000;
defparam ram16sdp_inst_465.INIT_2 = 16'h0000;
defparam ram16sdp_inst_465.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_466 (
    .DO(ram16sdp_inst_466_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_176),
    .CLK(clk)
);

defparam ram16sdp_inst_466.INIT_0 = 16'h0000;
defparam ram16sdp_inst_466.INIT_1 = 16'h0000;
defparam ram16sdp_inst_466.INIT_2 = 16'h0000;
defparam ram16sdp_inst_466.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_467 (
    .DO(ram16sdp_inst_467_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_176),
    .CLK(clk)
);

defparam ram16sdp_inst_467.INIT_0 = 16'h0000;
defparam ram16sdp_inst_467.INIT_1 = 16'h0000;
defparam ram16sdp_inst_467.INIT_2 = 16'h0000;
defparam ram16sdp_inst_467.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_468 (
    .DO(ram16sdp_inst_468_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_176),
    .CLK(clk)
);

defparam ram16sdp_inst_468.INIT_0 = 16'h0000;
defparam ram16sdp_inst_468.INIT_1 = 16'h0000;
defparam ram16sdp_inst_468.INIT_2 = 16'h0000;
defparam ram16sdp_inst_468.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_469 (
    .DO(ram16sdp_inst_469_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_176),
    .CLK(clk)
);

defparam ram16sdp_inst_469.INIT_0 = 16'h0000;
defparam ram16sdp_inst_469.INIT_1 = 16'h0000;
defparam ram16sdp_inst_469.INIT_2 = 16'h0000;
defparam ram16sdp_inst_469.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_470 (
    .DO(ram16sdp_inst_470_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_176),
    .CLK(clk)
);

defparam ram16sdp_inst_470.INIT_0 = 16'h0000;
defparam ram16sdp_inst_470.INIT_1 = 16'h0000;
defparam ram16sdp_inst_470.INIT_2 = 16'h0000;
defparam ram16sdp_inst_470.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_471 (
    .DO(ram16sdp_inst_471_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_176),
    .CLK(clk)
);

defparam ram16sdp_inst_471.INIT_0 = 16'h0000;
defparam ram16sdp_inst_471.INIT_1 = 16'h0000;
defparam ram16sdp_inst_471.INIT_2 = 16'h0000;
defparam ram16sdp_inst_471.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_472 (
    .DO(ram16sdp_inst_472_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16sdp_inst_472.INIT_0 = 16'h0000;
defparam ram16sdp_inst_472.INIT_1 = 16'h0000;
defparam ram16sdp_inst_472.INIT_2 = 16'h0000;
defparam ram16sdp_inst_472.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_473 (
    .DO(ram16sdp_inst_473_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16sdp_inst_473.INIT_0 = 16'h0000;
defparam ram16sdp_inst_473.INIT_1 = 16'h0000;
defparam ram16sdp_inst_473.INIT_2 = 16'h0000;
defparam ram16sdp_inst_473.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_474 (
    .DO(ram16sdp_inst_474_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16sdp_inst_474.INIT_0 = 16'h0000;
defparam ram16sdp_inst_474.INIT_1 = 16'h0000;
defparam ram16sdp_inst_474.INIT_2 = 16'h0000;
defparam ram16sdp_inst_474.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_475 (
    .DO(ram16sdp_inst_475_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16sdp_inst_475.INIT_0 = 16'h0000;
defparam ram16sdp_inst_475.INIT_1 = 16'h0000;
defparam ram16sdp_inst_475.INIT_2 = 16'h0000;
defparam ram16sdp_inst_475.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_476 (
    .DO(ram16sdp_inst_476_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16sdp_inst_476.INIT_0 = 16'h0000;
defparam ram16sdp_inst_476.INIT_1 = 16'h0000;
defparam ram16sdp_inst_476.INIT_2 = 16'h0000;
defparam ram16sdp_inst_476.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_477 (
    .DO(ram16sdp_inst_477_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16sdp_inst_477.INIT_0 = 16'h0000;
defparam ram16sdp_inst_477.INIT_1 = 16'h0000;
defparam ram16sdp_inst_477.INIT_2 = 16'h0000;
defparam ram16sdp_inst_477.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_478 (
    .DO(ram16sdp_inst_478_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16sdp_inst_478.INIT_0 = 16'h0000;
defparam ram16sdp_inst_478.INIT_1 = 16'h0000;
defparam ram16sdp_inst_478.INIT_2 = 16'h0000;
defparam ram16sdp_inst_478.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_479 (
    .DO(ram16sdp_inst_479_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16sdp_inst_479.INIT_0 = 16'h0000;
defparam ram16sdp_inst_479.INIT_1 = 16'h0000;
defparam ram16sdp_inst_479.INIT_2 = 16'h0000;
defparam ram16sdp_inst_479.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_480 (
    .DO(ram16sdp_inst_480_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_182),
    .CLK(clk)
);

defparam ram16sdp_inst_480.INIT_0 = 16'h0000;
defparam ram16sdp_inst_480.INIT_1 = 16'h0000;
defparam ram16sdp_inst_480.INIT_2 = 16'h0000;
defparam ram16sdp_inst_480.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_481 (
    .DO(ram16sdp_inst_481_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_182),
    .CLK(clk)
);

defparam ram16sdp_inst_481.INIT_0 = 16'h0000;
defparam ram16sdp_inst_481.INIT_1 = 16'h0000;
defparam ram16sdp_inst_481.INIT_2 = 16'h0000;
defparam ram16sdp_inst_481.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_482 (
    .DO(ram16sdp_inst_482_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_182),
    .CLK(clk)
);

defparam ram16sdp_inst_482.INIT_0 = 16'h0000;
defparam ram16sdp_inst_482.INIT_1 = 16'h0000;
defparam ram16sdp_inst_482.INIT_2 = 16'h0000;
defparam ram16sdp_inst_482.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_483 (
    .DO(ram16sdp_inst_483_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_182),
    .CLK(clk)
);

defparam ram16sdp_inst_483.INIT_0 = 16'h0000;
defparam ram16sdp_inst_483.INIT_1 = 16'h0000;
defparam ram16sdp_inst_483.INIT_2 = 16'h0000;
defparam ram16sdp_inst_483.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_484 (
    .DO(ram16sdp_inst_484_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_182),
    .CLK(clk)
);

defparam ram16sdp_inst_484.INIT_0 = 16'h0000;
defparam ram16sdp_inst_484.INIT_1 = 16'h0000;
defparam ram16sdp_inst_484.INIT_2 = 16'h0000;
defparam ram16sdp_inst_484.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_485 (
    .DO(ram16sdp_inst_485_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_182),
    .CLK(clk)
);

defparam ram16sdp_inst_485.INIT_0 = 16'h0000;
defparam ram16sdp_inst_485.INIT_1 = 16'h0000;
defparam ram16sdp_inst_485.INIT_2 = 16'h0000;
defparam ram16sdp_inst_485.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_486 (
    .DO(ram16sdp_inst_486_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_182),
    .CLK(clk)
);

defparam ram16sdp_inst_486.INIT_0 = 16'h0000;
defparam ram16sdp_inst_486.INIT_1 = 16'h0000;
defparam ram16sdp_inst_486.INIT_2 = 16'h0000;
defparam ram16sdp_inst_486.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_487 (
    .DO(ram16sdp_inst_487_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_182),
    .CLK(clk)
);

defparam ram16sdp_inst_487.INIT_0 = 16'h0000;
defparam ram16sdp_inst_487.INIT_1 = 16'h0000;
defparam ram16sdp_inst_487.INIT_2 = 16'h0000;
defparam ram16sdp_inst_487.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_488 (
    .DO(ram16sdp_inst_488_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_185),
    .CLK(clk)
);

defparam ram16sdp_inst_488.INIT_0 = 16'h0000;
defparam ram16sdp_inst_488.INIT_1 = 16'h0000;
defparam ram16sdp_inst_488.INIT_2 = 16'h0000;
defparam ram16sdp_inst_488.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_489 (
    .DO(ram16sdp_inst_489_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_185),
    .CLK(clk)
);

defparam ram16sdp_inst_489.INIT_0 = 16'h0000;
defparam ram16sdp_inst_489.INIT_1 = 16'h0000;
defparam ram16sdp_inst_489.INIT_2 = 16'h0000;
defparam ram16sdp_inst_489.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_490 (
    .DO(ram16sdp_inst_490_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_185),
    .CLK(clk)
);

defparam ram16sdp_inst_490.INIT_0 = 16'h0000;
defparam ram16sdp_inst_490.INIT_1 = 16'h0000;
defparam ram16sdp_inst_490.INIT_2 = 16'h0000;
defparam ram16sdp_inst_490.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_491 (
    .DO(ram16sdp_inst_491_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_185),
    .CLK(clk)
);

defparam ram16sdp_inst_491.INIT_0 = 16'h0000;
defparam ram16sdp_inst_491.INIT_1 = 16'h0000;
defparam ram16sdp_inst_491.INIT_2 = 16'h0000;
defparam ram16sdp_inst_491.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_492 (
    .DO(ram16sdp_inst_492_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_185),
    .CLK(clk)
);

defparam ram16sdp_inst_492.INIT_0 = 16'h0000;
defparam ram16sdp_inst_492.INIT_1 = 16'h0000;
defparam ram16sdp_inst_492.INIT_2 = 16'h0000;
defparam ram16sdp_inst_492.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_493 (
    .DO(ram16sdp_inst_493_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_185),
    .CLK(clk)
);

defparam ram16sdp_inst_493.INIT_0 = 16'h0000;
defparam ram16sdp_inst_493.INIT_1 = 16'h0000;
defparam ram16sdp_inst_493.INIT_2 = 16'h0000;
defparam ram16sdp_inst_493.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_494 (
    .DO(ram16sdp_inst_494_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_185),
    .CLK(clk)
);

defparam ram16sdp_inst_494.INIT_0 = 16'h0000;
defparam ram16sdp_inst_494.INIT_1 = 16'h0000;
defparam ram16sdp_inst_494.INIT_2 = 16'h0000;
defparam ram16sdp_inst_494.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_495 (
    .DO(ram16sdp_inst_495_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_185),
    .CLK(clk)
);

defparam ram16sdp_inst_495.INIT_0 = 16'h0000;
defparam ram16sdp_inst_495.INIT_1 = 16'h0000;
defparam ram16sdp_inst_495.INIT_2 = 16'h0000;
defparam ram16sdp_inst_495.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_496 (
    .DO(ram16sdp_inst_496_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_188),
    .CLK(clk)
);

defparam ram16sdp_inst_496.INIT_0 = 16'h0000;
defparam ram16sdp_inst_496.INIT_1 = 16'h0000;
defparam ram16sdp_inst_496.INIT_2 = 16'h0000;
defparam ram16sdp_inst_496.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_497 (
    .DO(ram16sdp_inst_497_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_188),
    .CLK(clk)
);

defparam ram16sdp_inst_497.INIT_0 = 16'h0000;
defparam ram16sdp_inst_497.INIT_1 = 16'h0000;
defparam ram16sdp_inst_497.INIT_2 = 16'h0000;
defparam ram16sdp_inst_497.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_498 (
    .DO(ram16sdp_inst_498_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_188),
    .CLK(clk)
);

defparam ram16sdp_inst_498.INIT_0 = 16'h0000;
defparam ram16sdp_inst_498.INIT_1 = 16'h0000;
defparam ram16sdp_inst_498.INIT_2 = 16'h0000;
defparam ram16sdp_inst_498.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_499 (
    .DO(ram16sdp_inst_499_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_188),
    .CLK(clk)
);

defparam ram16sdp_inst_499.INIT_0 = 16'h0000;
defparam ram16sdp_inst_499.INIT_1 = 16'h0000;
defparam ram16sdp_inst_499.INIT_2 = 16'h0000;
defparam ram16sdp_inst_499.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_500 (
    .DO(ram16sdp_inst_500_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_188),
    .CLK(clk)
);

defparam ram16sdp_inst_500.INIT_0 = 16'h0000;
defparam ram16sdp_inst_500.INIT_1 = 16'h0000;
defparam ram16sdp_inst_500.INIT_2 = 16'h0000;
defparam ram16sdp_inst_500.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_501 (
    .DO(ram16sdp_inst_501_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_188),
    .CLK(clk)
);

defparam ram16sdp_inst_501.INIT_0 = 16'h0000;
defparam ram16sdp_inst_501.INIT_1 = 16'h0000;
defparam ram16sdp_inst_501.INIT_2 = 16'h0000;
defparam ram16sdp_inst_501.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_502 (
    .DO(ram16sdp_inst_502_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_188),
    .CLK(clk)
);

defparam ram16sdp_inst_502.INIT_0 = 16'h0000;
defparam ram16sdp_inst_502.INIT_1 = 16'h0000;
defparam ram16sdp_inst_502.INIT_2 = 16'h0000;
defparam ram16sdp_inst_502.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_503 (
    .DO(ram16sdp_inst_503_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_188),
    .CLK(clk)
);

defparam ram16sdp_inst_503.INIT_0 = 16'h0000;
defparam ram16sdp_inst_503.INIT_1 = 16'h0000;
defparam ram16sdp_inst_503.INIT_2 = 16'h0000;
defparam ram16sdp_inst_503.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_504 (
    .DO(ram16sdp_inst_504_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16sdp_inst_504.INIT_0 = 16'h0000;
defparam ram16sdp_inst_504.INIT_1 = 16'h0000;
defparam ram16sdp_inst_504.INIT_2 = 16'h0000;
defparam ram16sdp_inst_504.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_505 (
    .DO(ram16sdp_inst_505_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16sdp_inst_505.INIT_0 = 16'h0000;
defparam ram16sdp_inst_505.INIT_1 = 16'h0000;
defparam ram16sdp_inst_505.INIT_2 = 16'h0000;
defparam ram16sdp_inst_505.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_506 (
    .DO(ram16sdp_inst_506_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16sdp_inst_506.INIT_0 = 16'h0000;
defparam ram16sdp_inst_506.INIT_1 = 16'h0000;
defparam ram16sdp_inst_506.INIT_2 = 16'h0000;
defparam ram16sdp_inst_506.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_507 (
    .DO(ram16sdp_inst_507_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16sdp_inst_507.INIT_0 = 16'h0000;
defparam ram16sdp_inst_507.INIT_1 = 16'h0000;
defparam ram16sdp_inst_507.INIT_2 = 16'h0000;
defparam ram16sdp_inst_507.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_508 (
    .DO(ram16sdp_inst_508_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16sdp_inst_508.INIT_0 = 16'h0000;
defparam ram16sdp_inst_508.INIT_1 = 16'h0000;
defparam ram16sdp_inst_508.INIT_2 = 16'h0000;
defparam ram16sdp_inst_508.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_509 (
    .DO(ram16sdp_inst_509_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16sdp_inst_509.INIT_0 = 16'h0000;
defparam ram16sdp_inst_509.INIT_1 = 16'h0000;
defparam ram16sdp_inst_509.INIT_2 = 16'h0000;
defparam ram16sdp_inst_509.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_510 (
    .DO(ram16sdp_inst_510_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16sdp_inst_510.INIT_0 = 16'h0000;
defparam ram16sdp_inst_510.INIT_1 = 16'h0000;
defparam ram16sdp_inst_510.INIT_2 = 16'h0000;
defparam ram16sdp_inst_510.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_511 (
    .DO(ram16sdp_inst_511_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16sdp_inst_511.INIT_0 = 16'h0000;
defparam ram16sdp_inst_511.INIT_1 = 16'h0000;
defparam ram16sdp_inst_511.INIT_2 = 16'h0000;
defparam ram16sdp_inst_511.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_512 (
    .DO(ram16sdp_inst_512_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_194),
    .CLK(clk)
);

defparam ram16sdp_inst_512.INIT_0 = 16'h0000;
defparam ram16sdp_inst_512.INIT_1 = 16'h0000;
defparam ram16sdp_inst_512.INIT_2 = 16'h0000;
defparam ram16sdp_inst_512.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_513 (
    .DO(ram16sdp_inst_513_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_194),
    .CLK(clk)
);

defparam ram16sdp_inst_513.INIT_0 = 16'h0000;
defparam ram16sdp_inst_513.INIT_1 = 16'h0000;
defparam ram16sdp_inst_513.INIT_2 = 16'h0000;
defparam ram16sdp_inst_513.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_514 (
    .DO(ram16sdp_inst_514_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_194),
    .CLK(clk)
);

defparam ram16sdp_inst_514.INIT_0 = 16'h0000;
defparam ram16sdp_inst_514.INIT_1 = 16'h0000;
defparam ram16sdp_inst_514.INIT_2 = 16'h0000;
defparam ram16sdp_inst_514.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_515 (
    .DO(ram16sdp_inst_515_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_194),
    .CLK(clk)
);

defparam ram16sdp_inst_515.INIT_0 = 16'h0000;
defparam ram16sdp_inst_515.INIT_1 = 16'h0000;
defparam ram16sdp_inst_515.INIT_2 = 16'h0000;
defparam ram16sdp_inst_515.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_516 (
    .DO(ram16sdp_inst_516_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_194),
    .CLK(clk)
);

defparam ram16sdp_inst_516.INIT_0 = 16'h0000;
defparam ram16sdp_inst_516.INIT_1 = 16'h0000;
defparam ram16sdp_inst_516.INIT_2 = 16'h0000;
defparam ram16sdp_inst_516.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_517 (
    .DO(ram16sdp_inst_517_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_194),
    .CLK(clk)
);

defparam ram16sdp_inst_517.INIT_0 = 16'h0000;
defparam ram16sdp_inst_517.INIT_1 = 16'h0000;
defparam ram16sdp_inst_517.INIT_2 = 16'h0000;
defparam ram16sdp_inst_517.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_518 (
    .DO(ram16sdp_inst_518_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_194),
    .CLK(clk)
);

defparam ram16sdp_inst_518.INIT_0 = 16'h0000;
defparam ram16sdp_inst_518.INIT_1 = 16'h0000;
defparam ram16sdp_inst_518.INIT_2 = 16'h0000;
defparam ram16sdp_inst_518.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_519 (
    .DO(ram16sdp_inst_519_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_194),
    .CLK(clk)
);

defparam ram16sdp_inst_519.INIT_0 = 16'h0000;
defparam ram16sdp_inst_519.INIT_1 = 16'h0000;
defparam ram16sdp_inst_519.INIT_2 = 16'h0000;
defparam ram16sdp_inst_519.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_520 (
    .DO(ram16sdp_inst_520_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_197),
    .CLK(clk)
);

defparam ram16sdp_inst_520.INIT_0 = 16'h0000;
defparam ram16sdp_inst_520.INIT_1 = 16'h0000;
defparam ram16sdp_inst_520.INIT_2 = 16'h0000;
defparam ram16sdp_inst_520.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_521 (
    .DO(ram16sdp_inst_521_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_197),
    .CLK(clk)
);

defparam ram16sdp_inst_521.INIT_0 = 16'h0000;
defparam ram16sdp_inst_521.INIT_1 = 16'h0000;
defparam ram16sdp_inst_521.INIT_2 = 16'h0000;
defparam ram16sdp_inst_521.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_522 (
    .DO(ram16sdp_inst_522_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_197),
    .CLK(clk)
);

defparam ram16sdp_inst_522.INIT_0 = 16'h0000;
defparam ram16sdp_inst_522.INIT_1 = 16'h0000;
defparam ram16sdp_inst_522.INIT_2 = 16'h0000;
defparam ram16sdp_inst_522.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_523 (
    .DO(ram16sdp_inst_523_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_197),
    .CLK(clk)
);

defparam ram16sdp_inst_523.INIT_0 = 16'h0000;
defparam ram16sdp_inst_523.INIT_1 = 16'h0000;
defparam ram16sdp_inst_523.INIT_2 = 16'h0000;
defparam ram16sdp_inst_523.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_524 (
    .DO(ram16sdp_inst_524_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_197),
    .CLK(clk)
);

defparam ram16sdp_inst_524.INIT_0 = 16'h0000;
defparam ram16sdp_inst_524.INIT_1 = 16'h0000;
defparam ram16sdp_inst_524.INIT_2 = 16'h0000;
defparam ram16sdp_inst_524.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_525 (
    .DO(ram16sdp_inst_525_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_197),
    .CLK(clk)
);

defparam ram16sdp_inst_525.INIT_0 = 16'h0000;
defparam ram16sdp_inst_525.INIT_1 = 16'h0000;
defparam ram16sdp_inst_525.INIT_2 = 16'h0000;
defparam ram16sdp_inst_525.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_526 (
    .DO(ram16sdp_inst_526_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_197),
    .CLK(clk)
);

defparam ram16sdp_inst_526.INIT_0 = 16'h0000;
defparam ram16sdp_inst_526.INIT_1 = 16'h0000;
defparam ram16sdp_inst_526.INIT_2 = 16'h0000;
defparam ram16sdp_inst_526.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_527 (
    .DO(ram16sdp_inst_527_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_197),
    .CLK(clk)
);

defparam ram16sdp_inst_527.INIT_0 = 16'h0000;
defparam ram16sdp_inst_527.INIT_1 = 16'h0000;
defparam ram16sdp_inst_527.INIT_2 = 16'h0000;
defparam ram16sdp_inst_527.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_528 (
    .DO(ram16sdp_inst_528_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_200),
    .CLK(clk)
);

defparam ram16sdp_inst_528.INIT_0 = 16'h0000;
defparam ram16sdp_inst_528.INIT_1 = 16'h0000;
defparam ram16sdp_inst_528.INIT_2 = 16'h0000;
defparam ram16sdp_inst_528.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_529 (
    .DO(ram16sdp_inst_529_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_200),
    .CLK(clk)
);

defparam ram16sdp_inst_529.INIT_0 = 16'h0000;
defparam ram16sdp_inst_529.INIT_1 = 16'h0000;
defparam ram16sdp_inst_529.INIT_2 = 16'h0000;
defparam ram16sdp_inst_529.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_530 (
    .DO(ram16sdp_inst_530_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_200),
    .CLK(clk)
);

defparam ram16sdp_inst_530.INIT_0 = 16'h0000;
defparam ram16sdp_inst_530.INIT_1 = 16'h0000;
defparam ram16sdp_inst_530.INIT_2 = 16'h0000;
defparam ram16sdp_inst_530.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_531 (
    .DO(ram16sdp_inst_531_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_200),
    .CLK(clk)
);

defparam ram16sdp_inst_531.INIT_0 = 16'h0000;
defparam ram16sdp_inst_531.INIT_1 = 16'h0000;
defparam ram16sdp_inst_531.INIT_2 = 16'h0000;
defparam ram16sdp_inst_531.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_532 (
    .DO(ram16sdp_inst_532_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_200),
    .CLK(clk)
);

defparam ram16sdp_inst_532.INIT_0 = 16'h0000;
defparam ram16sdp_inst_532.INIT_1 = 16'h0000;
defparam ram16sdp_inst_532.INIT_2 = 16'h0000;
defparam ram16sdp_inst_532.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_533 (
    .DO(ram16sdp_inst_533_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_200),
    .CLK(clk)
);

defparam ram16sdp_inst_533.INIT_0 = 16'h0000;
defparam ram16sdp_inst_533.INIT_1 = 16'h0000;
defparam ram16sdp_inst_533.INIT_2 = 16'h0000;
defparam ram16sdp_inst_533.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_534 (
    .DO(ram16sdp_inst_534_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_200),
    .CLK(clk)
);

defparam ram16sdp_inst_534.INIT_0 = 16'h0000;
defparam ram16sdp_inst_534.INIT_1 = 16'h0000;
defparam ram16sdp_inst_534.INIT_2 = 16'h0000;
defparam ram16sdp_inst_534.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_535 (
    .DO(ram16sdp_inst_535_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_200),
    .CLK(clk)
);

defparam ram16sdp_inst_535.INIT_0 = 16'h0000;
defparam ram16sdp_inst_535.INIT_1 = 16'h0000;
defparam ram16sdp_inst_535.INIT_2 = 16'h0000;
defparam ram16sdp_inst_535.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_536 (
    .DO(ram16sdp_inst_536_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16sdp_inst_536.INIT_0 = 16'h0000;
defparam ram16sdp_inst_536.INIT_1 = 16'h0000;
defparam ram16sdp_inst_536.INIT_2 = 16'h0000;
defparam ram16sdp_inst_536.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_537 (
    .DO(ram16sdp_inst_537_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16sdp_inst_537.INIT_0 = 16'h0000;
defparam ram16sdp_inst_537.INIT_1 = 16'h0000;
defparam ram16sdp_inst_537.INIT_2 = 16'h0000;
defparam ram16sdp_inst_537.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_538 (
    .DO(ram16sdp_inst_538_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16sdp_inst_538.INIT_0 = 16'h0000;
defparam ram16sdp_inst_538.INIT_1 = 16'h0000;
defparam ram16sdp_inst_538.INIT_2 = 16'h0000;
defparam ram16sdp_inst_538.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_539 (
    .DO(ram16sdp_inst_539_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16sdp_inst_539.INIT_0 = 16'h0000;
defparam ram16sdp_inst_539.INIT_1 = 16'h0000;
defparam ram16sdp_inst_539.INIT_2 = 16'h0000;
defparam ram16sdp_inst_539.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_540 (
    .DO(ram16sdp_inst_540_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16sdp_inst_540.INIT_0 = 16'h0000;
defparam ram16sdp_inst_540.INIT_1 = 16'h0000;
defparam ram16sdp_inst_540.INIT_2 = 16'h0000;
defparam ram16sdp_inst_540.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_541 (
    .DO(ram16sdp_inst_541_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16sdp_inst_541.INIT_0 = 16'h0000;
defparam ram16sdp_inst_541.INIT_1 = 16'h0000;
defparam ram16sdp_inst_541.INIT_2 = 16'h0000;
defparam ram16sdp_inst_541.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_542 (
    .DO(ram16sdp_inst_542_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16sdp_inst_542.INIT_0 = 16'h0000;
defparam ram16sdp_inst_542.INIT_1 = 16'h0000;
defparam ram16sdp_inst_542.INIT_2 = 16'h0000;
defparam ram16sdp_inst_542.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_543 (
    .DO(ram16sdp_inst_543_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16sdp_inst_543.INIT_0 = 16'h0000;
defparam ram16sdp_inst_543.INIT_1 = 16'h0000;
defparam ram16sdp_inst_543.INIT_2 = 16'h0000;
defparam ram16sdp_inst_543.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_544 (
    .DO(ram16sdp_inst_544_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_206),
    .CLK(clk)
);

defparam ram16sdp_inst_544.INIT_0 = 16'h0000;
defparam ram16sdp_inst_544.INIT_1 = 16'h0000;
defparam ram16sdp_inst_544.INIT_2 = 16'h0000;
defparam ram16sdp_inst_544.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_545 (
    .DO(ram16sdp_inst_545_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_206),
    .CLK(clk)
);

defparam ram16sdp_inst_545.INIT_0 = 16'h0000;
defparam ram16sdp_inst_545.INIT_1 = 16'h0000;
defparam ram16sdp_inst_545.INIT_2 = 16'h0000;
defparam ram16sdp_inst_545.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_546 (
    .DO(ram16sdp_inst_546_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_206),
    .CLK(clk)
);

defparam ram16sdp_inst_546.INIT_0 = 16'h0000;
defparam ram16sdp_inst_546.INIT_1 = 16'h0000;
defparam ram16sdp_inst_546.INIT_2 = 16'h0000;
defparam ram16sdp_inst_546.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_547 (
    .DO(ram16sdp_inst_547_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_206),
    .CLK(clk)
);

defparam ram16sdp_inst_547.INIT_0 = 16'h0000;
defparam ram16sdp_inst_547.INIT_1 = 16'h0000;
defparam ram16sdp_inst_547.INIT_2 = 16'h0000;
defparam ram16sdp_inst_547.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_548 (
    .DO(ram16sdp_inst_548_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_206),
    .CLK(clk)
);

defparam ram16sdp_inst_548.INIT_0 = 16'h0000;
defparam ram16sdp_inst_548.INIT_1 = 16'h0000;
defparam ram16sdp_inst_548.INIT_2 = 16'h0000;
defparam ram16sdp_inst_548.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_549 (
    .DO(ram16sdp_inst_549_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_206),
    .CLK(clk)
);

defparam ram16sdp_inst_549.INIT_0 = 16'h0000;
defparam ram16sdp_inst_549.INIT_1 = 16'h0000;
defparam ram16sdp_inst_549.INIT_2 = 16'h0000;
defparam ram16sdp_inst_549.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_550 (
    .DO(ram16sdp_inst_550_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_206),
    .CLK(clk)
);

defparam ram16sdp_inst_550.INIT_0 = 16'h0000;
defparam ram16sdp_inst_550.INIT_1 = 16'h0000;
defparam ram16sdp_inst_550.INIT_2 = 16'h0000;
defparam ram16sdp_inst_550.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_551 (
    .DO(ram16sdp_inst_551_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_206),
    .CLK(clk)
);

defparam ram16sdp_inst_551.INIT_0 = 16'h0000;
defparam ram16sdp_inst_551.INIT_1 = 16'h0000;
defparam ram16sdp_inst_551.INIT_2 = 16'h0000;
defparam ram16sdp_inst_551.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_552 (
    .DO(ram16sdp_inst_552_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_209),
    .CLK(clk)
);

defparam ram16sdp_inst_552.INIT_0 = 16'h0000;
defparam ram16sdp_inst_552.INIT_1 = 16'h0000;
defparam ram16sdp_inst_552.INIT_2 = 16'h0000;
defparam ram16sdp_inst_552.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_553 (
    .DO(ram16sdp_inst_553_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_209),
    .CLK(clk)
);

defparam ram16sdp_inst_553.INIT_0 = 16'h0000;
defparam ram16sdp_inst_553.INIT_1 = 16'h0000;
defparam ram16sdp_inst_553.INIT_2 = 16'h0000;
defparam ram16sdp_inst_553.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_554 (
    .DO(ram16sdp_inst_554_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_209),
    .CLK(clk)
);

defparam ram16sdp_inst_554.INIT_0 = 16'h0000;
defparam ram16sdp_inst_554.INIT_1 = 16'h0000;
defparam ram16sdp_inst_554.INIT_2 = 16'h0000;
defparam ram16sdp_inst_554.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_555 (
    .DO(ram16sdp_inst_555_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_209),
    .CLK(clk)
);

defparam ram16sdp_inst_555.INIT_0 = 16'h0000;
defparam ram16sdp_inst_555.INIT_1 = 16'h0000;
defparam ram16sdp_inst_555.INIT_2 = 16'h0000;
defparam ram16sdp_inst_555.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_556 (
    .DO(ram16sdp_inst_556_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_209),
    .CLK(clk)
);

defparam ram16sdp_inst_556.INIT_0 = 16'h0000;
defparam ram16sdp_inst_556.INIT_1 = 16'h0000;
defparam ram16sdp_inst_556.INIT_2 = 16'h0000;
defparam ram16sdp_inst_556.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_557 (
    .DO(ram16sdp_inst_557_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_209),
    .CLK(clk)
);

defparam ram16sdp_inst_557.INIT_0 = 16'h0000;
defparam ram16sdp_inst_557.INIT_1 = 16'h0000;
defparam ram16sdp_inst_557.INIT_2 = 16'h0000;
defparam ram16sdp_inst_557.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_558 (
    .DO(ram16sdp_inst_558_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_209),
    .CLK(clk)
);

defparam ram16sdp_inst_558.INIT_0 = 16'h0000;
defparam ram16sdp_inst_558.INIT_1 = 16'h0000;
defparam ram16sdp_inst_558.INIT_2 = 16'h0000;
defparam ram16sdp_inst_558.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_559 (
    .DO(ram16sdp_inst_559_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_209),
    .CLK(clk)
);

defparam ram16sdp_inst_559.INIT_0 = 16'h0000;
defparam ram16sdp_inst_559.INIT_1 = 16'h0000;
defparam ram16sdp_inst_559.INIT_2 = 16'h0000;
defparam ram16sdp_inst_559.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_560 (
    .DO(ram16sdp_inst_560_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_212),
    .CLK(clk)
);

defparam ram16sdp_inst_560.INIT_0 = 16'h0000;
defparam ram16sdp_inst_560.INIT_1 = 16'h0000;
defparam ram16sdp_inst_560.INIT_2 = 16'h0000;
defparam ram16sdp_inst_560.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_561 (
    .DO(ram16sdp_inst_561_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_212),
    .CLK(clk)
);

defparam ram16sdp_inst_561.INIT_0 = 16'h0000;
defparam ram16sdp_inst_561.INIT_1 = 16'h0000;
defparam ram16sdp_inst_561.INIT_2 = 16'h0000;
defparam ram16sdp_inst_561.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_562 (
    .DO(ram16sdp_inst_562_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_212),
    .CLK(clk)
);

defparam ram16sdp_inst_562.INIT_0 = 16'h0000;
defparam ram16sdp_inst_562.INIT_1 = 16'h0000;
defparam ram16sdp_inst_562.INIT_2 = 16'h0000;
defparam ram16sdp_inst_562.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_563 (
    .DO(ram16sdp_inst_563_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_212),
    .CLK(clk)
);

defparam ram16sdp_inst_563.INIT_0 = 16'h0000;
defparam ram16sdp_inst_563.INIT_1 = 16'h0000;
defparam ram16sdp_inst_563.INIT_2 = 16'h0000;
defparam ram16sdp_inst_563.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_564 (
    .DO(ram16sdp_inst_564_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_212),
    .CLK(clk)
);

defparam ram16sdp_inst_564.INIT_0 = 16'h0000;
defparam ram16sdp_inst_564.INIT_1 = 16'h0000;
defparam ram16sdp_inst_564.INIT_2 = 16'h0000;
defparam ram16sdp_inst_564.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_565 (
    .DO(ram16sdp_inst_565_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_212),
    .CLK(clk)
);

defparam ram16sdp_inst_565.INIT_0 = 16'h0000;
defparam ram16sdp_inst_565.INIT_1 = 16'h0000;
defparam ram16sdp_inst_565.INIT_2 = 16'h0000;
defparam ram16sdp_inst_565.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_566 (
    .DO(ram16sdp_inst_566_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_212),
    .CLK(clk)
);

defparam ram16sdp_inst_566.INIT_0 = 16'h0000;
defparam ram16sdp_inst_566.INIT_1 = 16'h0000;
defparam ram16sdp_inst_566.INIT_2 = 16'h0000;
defparam ram16sdp_inst_566.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_567 (
    .DO(ram16sdp_inst_567_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_212),
    .CLK(clk)
);

defparam ram16sdp_inst_567.INIT_0 = 16'h0000;
defparam ram16sdp_inst_567.INIT_1 = 16'h0000;
defparam ram16sdp_inst_567.INIT_2 = 16'h0000;
defparam ram16sdp_inst_567.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_568 (
    .DO(ram16sdp_inst_568_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16sdp_inst_568.INIT_0 = 16'h0000;
defparam ram16sdp_inst_568.INIT_1 = 16'h0000;
defparam ram16sdp_inst_568.INIT_2 = 16'h0000;
defparam ram16sdp_inst_568.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_569 (
    .DO(ram16sdp_inst_569_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16sdp_inst_569.INIT_0 = 16'h0000;
defparam ram16sdp_inst_569.INIT_1 = 16'h0000;
defparam ram16sdp_inst_569.INIT_2 = 16'h0000;
defparam ram16sdp_inst_569.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_570 (
    .DO(ram16sdp_inst_570_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16sdp_inst_570.INIT_0 = 16'h0000;
defparam ram16sdp_inst_570.INIT_1 = 16'h0000;
defparam ram16sdp_inst_570.INIT_2 = 16'h0000;
defparam ram16sdp_inst_570.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_571 (
    .DO(ram16sdp_inst_571_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16sdp_inst_571.INIT_0 = 16'h0000;
defparam ram16sdp_inst_571.INIT_1 = 16'h0000;
defparam ram16sdp_inst_571.INIT_2 = 16'h0000;
defparam ram16sdp_inst_571.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_572 (
    .DO(ram16sdp_inst_572_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16sdp_inst_572.INIT_0 = 16'h0000;
defparam ram16sdp_inst_572.INIT_1 = 16'h0000;
defparam ram16sdp_inst_572.INIT_2 = 16'h0000;
defparam ram16sdp_inst_572.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_573 (
    .DO(ram16sdp_inst_573_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16sdp_inst_573.INIT_0 = 16'h0000;
defparam ram16sdp_inst_573.INIT_1 = 16'h0000;
defparam ram16sdp_inst_573.INIT_2 = 16'h0000;
defparam ram16sdp_inst_573.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_574 (
    .DO(ram16sdp_inst_574_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16sdp_inst_574.INIT_0 = 16'h0000;
defparam ram16sdp_inst_574.INIT_1 = 16'h0000;
defparam ram16sdp_inst_574.INIT_2 = 16'h0000;
defparam ram16sdp_inst_574.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_575 (
    .DO(ram16sdp_inst_575_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16sdp_inst_575.INIT_0 = 16'h0000;
defparam ram16sdp_inst_575.INIT_1 = 16'h0000;
defparam ram16sdp_inst_575.INIT_2 = 16'h0000;
defparam ram16sdp_inst_575.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_576 (
    .DO(ram16sdp_inst_576_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_218),
    .CLK(clk)
);

defparam ram16sdp_inst_576.INIT_0 = 16'h0000;
defparam ram16sdp_inst_576.INIT_1 = 16'h0000;
defparam ram16sdp_inst_576.INIT_2 = 16'h0000;
defparam ram16sdp_inst_576.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_577 (
    .DO(ram16sdp_inst_577_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_218),
    .CLK(clk)
);

defparam ram16sdp_inst_577.INIT_0 = 16'h0000;
defparam ram16sdp_inst_577.INIT_1 = 16'h0000;
defparam ram16sdp_inst_577.INIT_2 = 16'h0000;
defparam ram16sdp_inst_577.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_578 (
    .DO(ram16sdp_inst_578_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_218),
    .CLK(clk)
);

defparam ram16sdp_inst_578.INIT_0 = 16'h0000;
defparam ram16sdp_inst_578.INIT_1 = 16'h0000;
defparam ram16sdp_inst_578.INIT_2 = 16'h0000;
defparam ram16sdp_inst_578.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_579 (
    .DO(ram16sdp_inst_579_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_218),
    .CLK(clk)
);

defparam ram16sdp_inst_579.INIT_0 = 16'h0000;
defparam ram16sdp_inst_579.INIT_1 = 16'h0000;
defparam ram16sdp_inst_579.INIT_2 = 16'h0000;
defparam ram16sdp_inst_579.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_580 (
    .DO(ram16sdp_inst_580_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_218),
    .CLK(clk)
);

defparam ram16sdp_inst_580.INIT_0 = 16'h0000;
defparam ram16sdp_inst_580.INIT_1 = 16'h0000;
defparam ram16sdp_inst_580.INIT_2 = 16'h0000;
defparam ram16sdp_inst_580.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_581 (
    .DO(ram16sdp_inst_581_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_218),
    .CLK(clk)
);

defparam ram16sdp_inst_581.INIT_0 = 16'h0000;
defparam ram16sdp_inst_581.INIT_1 = 16'h0000;
defparam ram16sdp_inst_581.INIT_2 = 16'h0000;
defparam ram16sdp_inst_581.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_582 (
    .DO(ram16sdp_inst_582_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_218),
    .CLK(clk)
);

defparam ram16sdp_inst_582.INIT_0 = 16'h0000;
defparam ram16sdp_inst_582.INIT_1 = 16'h0000;
defparam ram16sdp_inst_582.INIT_2 = 16'h0000;
defparam ram16sdp_inst_582.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_583 (
    .DO(ram16sdp_inst_583_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_218),
    .CLK(clk)
);

defparam ram16sdp_inst_583.INIT_0 = 16'h0000;
defparam ram16sdp_inst_583.INIT_1 = 16'h0000;
defparam ram16sdp_inst_583.INIT_2 = 16'h0000;
defparam ram16sdp_inst_583.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_584 (
    .DO(ram16sdp_inst_584_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_221),
    .CLK(clk)
);

defparam ram16sdp_inst_584.INIT_0 = 16'h0000;
defparam ram16sdp_inst_584.INIT_1 = 16'h0000;
defparam ram16sdp_inst_584.INIT_2 = 16'h0000;
defparam ram16sdp_inst_584.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_585 (
    .DO(ram16sdp_inst_585_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_221),
    .CLK(clk)
);

defparam ram16sdp_inst_585.INIT_0 = 16'h0000;
defparam ram16sdp_inst_585.INIT_1 = 16'h0000;
defparam ram16sdp_inst_585.INIT_2 = 16'h0000;
defparam ram16sdp_inst_585.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_586 (
    .DO(ram16sdp_inst_586_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_221),
    .CLK(clk)
);

defparam ram16sdp_inst_586.INIT_0 = 16'h0000;
defparam ram16sdp_inst_586.INIT_1 = 16'h0000;
defparam ram16sdp_inst_586.INIT_2 = 16'h0000;
defparam ram16sdp_inst_586.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_587 (
    .DO(ram16sdp_inst_587_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_221),
    .CLK(clk)
);

defparam ram16sdp_inst_587.INIT_0 = 16'h0000;
defparam ram16sdp_inst_587.INIT_1 = 16'h0000;
defparam ram16sdp_inst_587.INIT_2 = 16'h0000;
defparam ram16sdp_inst_587.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_588 (
    .DO(ram16sdp_inst_588_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_221),
    .CLK(clk)
);

defparam ram16sdp_inst_588.INIT_0 = 16'h0000;
defparam ram16sdp_inst_588.INIT_1 = 16'h0000;
defparam ram16sdp_inst_588.INIT_2 = 16'h0000;
defparam ram16sdp_inst_588.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_589 (
    .DO(ram16sdp_inst_589_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_221),
    .CLK(clk)
);

defparam ram16sdp_inst_589.INIT_0 = 16'h0000;
defparam ram16sdp_inst_589.INIT_1 = 16'h0000;
defparam ram16sdp_inst_589.INIT_2 = 16'h0000;
defparam ram16sdp_inst_589.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_590 (
    .DO(ram16sdp_inst_590_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_221),
    .CLK(clk)
);

defparam ram16sdp_inst_590.INIT_0 = 16'h0000;
defparam ram16sdp_inst_590.INIT_1 = 16'h0000;
defparam ram16sdp_inst_590.INIT_2 = 16'h0000;
defparam ram16sdp_inst_590.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_591 (
    .DO(ram16sdp_inst_591_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_221),
    .CLK(clk)
);

defparam ram16sdp_inst_591.INIT_0 = 16'h0000;
defparam ram16sdp_inst_591.INIT_1 = 16'h0000;
defparam ram16sdp_inst_591.INIT_2 = 16'h0000;
defparam ram16sdp_inst_591.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_592 (
    .DO(ram16sdp_inst_592_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_224),
    .CLK(clk)
);

defparam ram16sdp_inst_592.INIT_0 = 16'h0000;
defparam ram16sdp_inst_592.INIT_1 = 16'h0000;
defparam ram16sdp_inst_592.INIT_2 = 16'h0000;
defparam ram16sdp_inst_592.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_593 (
    .DO(ram16sdp_inst_593_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_224),
    .CLK(clk)
);

defparam ram16sdp_inst_593.INIT_0 = 16'h0000;
defparam ram16sdp_inst_593.INIT_1 = 16'h0000;
defparam ram16sdp_inst_593.INIT_2 = 16'h0000;
defparam ram16sdp_inst_593.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_594 (
    .DO(ram16sdp_inst_594_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_224),
    .CLK(clk)
);

defparam ram16sdp_inst_594.INIT_0 = 16'h0000;
defparam ram16sdp_inst_594.INIT_1 = 16'h0000;
defparam ram16sdp_inst_594.INIT_2 = 16'h0000;
defparam ram16sdp_inst_594.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_595 (
    .DO(ram16sdp_inst_595_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_224),
    .CLK(clk)
);

defparam ram16sdp_inst_595.INIT_0 = 16'h0000;
defparam ram16sdp_inst_595.INIT_1 = 16'h0000;
defparam ram16sdp_inst_595.INIT_2 = 16'h0000;
defparam ram16sdp_inst_595.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_596 (
    .DO(ram16sdp_inst_596_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_224),
    .CLK(clk)
);

defparam ram16sdp_inst_596.INIT_0 = 16'h0000;
defparam ram16sdp_inst_596.INIT_1 = 16'h0000;
defparam ram16sdp_inst_596.INIT_2 = 16'h0000;
defparam ram16sdp_inst_596.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_597 (
    .DO(ram16sdp_inst_597_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_224),
    .CLK(clk)
);

defparam ram16sdp_inst_597.INIT_0 = 16'h0000;
defparam ram16sdp_inst_597.INIT_1 = 16'h0000;
defparam ram16sdp_inst_597.INIT_2 = 16'h0000;
defparam ram16sdp_inst_597.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_598 (
    .DO(ram16sdp_inst_598_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_224),
    .CLK(clk)
);

defparam ram16sdp_inst_598.INIT_0 = 16'h0000;
defparam ram16sdp_inst_598.INIT_1 = 16'h0000;
defparam ram16sdp_inst_598.INIT_2 = 16'h0000;
defparam ram16sdp_inst_598.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_599 (
    .DO(ram16sdp_inst_599_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_224),
    .CLK(clk)
);

defparam ram16sdp_inst_599.INIT_0 = 16'h0000;
defparam ram16sdp_inst_599.INIT_1 = 16'h0000;
defparam ram16sdp_inst_599.INIT_2 = 16'h0000;
defparam ram16sdp_inst_599.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_600 (
    .DO(ram16sdp_inst_600_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16sdp_inst_600.INIT_0 = 16'h0000;
defparam ram16sdp_inst_600.INIT_1 = 16'h0000;
defparam ram16sdp_inst_600.INIT_2 = 16'h0000;
defparam ram16sdp_inst_600.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_601 (
    .DO(ram16sdp_inst_601_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16sdp_inst_601.INIT_0 = 16'h0000;
defparam ram16sdp_inst_601.INIT_1 = 16'h0000;
defparam ram16sdp_inst_601.INIT_2 = 16'h0000;
defparam ram16sdp_inst_601.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_602 (
    .DO(ram16sdp_inst_602_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16sdp_inst_602.INIT_0 = 16'h0000;
defparam ram16sdp_inst_602.INIT_1 = 16'h0000;
defparam ram16sdp_inst_602.INIT_2 = 16'h0000;
defparam ram16sdp_inst_602.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_603 (
    .DO(ram16sdp_inst_603_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16sdp_inst_603.INIT_0 = 16'h0000;
defparam ram16sdp_inst_603.INIT_1 = 16'h0000;
defparam ram16sdp_inst_603.INIT_2 = 16'h0000;
defparam ram16sdp_inst_603.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_604 (
    .DO(ram16sdp_inst_604_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16sdp_inst_604.INIT_0 = 16'h0000;
defparam ram16sdp_inst_604.INIT_1 = 16'h0000;
defparam ram16sdp_inst_604.INIT_2 = 16'h0000;
defparam ram16sdp_inst_604.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_605 (
    .DO(ram16sdp_inst_605_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16sdp_inst_605.INIT_0 = 16'h0000;
defparam ram16sdp_inst_605.INIT_1 = 16'h0000;
defparam ram16sdp_inst_605.INIT_2 = 16'h0000;
defparam ram16sdp_inst_605.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_606 (
    .DO(ram16sdp_inst_606_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16sdp_inst_606.INIT_0 = 16'h0000;
defparam ram16sdp_inst_606.INIT_1 = 16'h0000;
defparam ram16sdp_inst_606.INIT_2 = 16'h0000;
defparam ram16sdp_inst_606.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_607 (
    .DO(ram16sdp_inst_607_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16sdp_inst_607.INIT_0 = 16'h0000;
defparam ram16sdp_inst_607.INIT_1 = 16'h0000;
defparam ram16sdp_inst_607.INIT_2 = 16'h0000;
defparam ram16sdp_inst_607.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_608 (
    .DO(ram16sdp_inst_608_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_230),
    .CLK(clk)
);

defparam ram16sdp_inst_608.INIT_0 = 16'h0000;
defparam ram16sdp_inst_608.INIT_1 = 16'h0000;
defparam ram16sdp_inst_608.INIT_2 = 16'h0000;
defparam ram16sdp_inst_608.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_609 (
    .DO(ram16sdp_inst_609_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_230),
    .CLK(clk)
);

defparam ram16sdp_inst_609.INIT_0 = 16'h0000;
defparam ram16sdp_inst_609.INIT_1 = 16'h0000;
defparam ram16sdp_inst_609.INIT_2 = 16'h0000;
defparam ram16sdp_inst_609.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_610 (
    .DO(ram16sdp_inst_610_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_230),
    .CLK(clk)
);

defparam ram16sdp_inst_610.INIT_0 = 16'h0000;
defparam ram16sdp_inst_610.INIT_1 = 16'h0000;
defparam ram16sdp_inst_610.INIT_2 = 16'h0000;
defparam ram16sdp_inst_610.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_611 (
    .DO(ram16sdp_inst_611_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_230),
    .CLK(clk)
);

defparam ram16sdp_inst_611.INIT_0 = 16'h0000;
defparam ram16sdp_inst_611.INIT_1 = 16'h0000;
defparam ram16sdp_inst_611.INIT_2 = 16'h0000;
defparam ram16sdp_inst_611.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_612 (
    .DO(ram16sdp_inst_612_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_230),
    .CLK(clk)
);

defparam ram16sdp_inst_612.INIT_0 = 16'h0000;
defparam ram16sdp_inst_612.INIT_1 = 16'h0000;
defparam ram16sdp_inst_612.INIT_2 = 16'h0000;
defparam ram16sdp_inst_612.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_613 (
    .DO(ram16sdp_inst_613_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_230),
    .CLK(clk)
);

defparam ram16sdp_inst_613.INIT_0 = 16'h0000;
defparam ram16sdp_inst_613.INIT_1 = 16'h0000;
defparam ram16sdp_inst_613.INIT_2 = 16'h0000;
defparam ram16sdp_inst_613.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_614 (
    .DO(ram16sdp_inst_614_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_230),
    .CLK(clk)
);

defparam ram16sdp_inst_614.INIT_0 = 16'h0000;
defparam ram16sdp_inst_614.INIT_1 = 16'h0000;
defparam ram16sdp_inst_614.INIT_2 = 16'h0000;
defparam ram16sdp_inst_614.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_615 (
    .DO(ram16sdp_inst_615_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_230),
    .CLK(clk)
);

defparam ram16sdp_inst_615.INIT_0 = 16'h0000;
defparam ram16sdp_inst_615.INIT_1 = 16'h0000;
defparam ram16sdp_inst_615.INIT_2 = 16'h0000;
defparam ram16sdp_inst_615.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_616 (
    .DO(ram16sdp_inst_616_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_233),
    .CLK(clk)
);

defparam ram16sdp_inst_616.INIT_0 = 16'h0000;
defparam ram16sdp_inst_616.INIT_1 = 16'h0000;
defparam ram16sdp_inst_616.INIT_2 = 16'h0000;
defparam ram16sdp_inst_616.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_617 (
    .DO(ram16sdp_inst_617_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_233),
    .CLK(clk)
);

defparam ram16sdp_inst_617.INIT_0 = 16'h0000;
defparam ram16sdp_inst_617.INIT_1 = 16'h0000;
defparam ram16sdp_inst_617.INIT_2 = 16'h0000;
defparam ram16sdp_inst_617.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_618 (
    .DO(ram16sdp_inst_618_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_233),
    .CLK(clk)
);

defparam ram16sdp_inst_618.INIT_0 = 16'h0000;
defparam ram16sdp_inst_618.INIT_1 = 16'h0000;
defparam ram16sdp_inst_618.INIT_2 = 16'h0000;
defparam ram16sdp_inst_618.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_619 (
    .DO(ram16sdp_inst_619_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_233),
    .CLK(clk)
);

defparam ram16sdp_inst_619.INIT_0 = 16'h0000;
defparam ram16sdp_inst_619.INIT_1 = 16'h0000;
defparam ram16sdp_inst_619.INIT_2 = 16'h0000;
defparam ram16sdp_inst_619.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_620 (
    .DO(ram16sdp_inst_620_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_233),
    .CLK(clk)
);

defparam ram16sdp_inst_620.INIT_0 = 16'h0000;
defparam ram16sdp_inst_620.INIT_1 = 16'h0000;
defparam ram16sdp_inst_620.INIT_2 = 16'h0000;
defparam ram16sdp_inst_620.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_621 (
    .DO(ram16sdp_inst_621_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_233),
    .CLK(clk)
);

defparam ram16sdp_inst_621.INIT_0 = 16'h0000;
defparam ram16sdp_inst_621.INIT_1 = 16'h0000;
defparam ram16sdp_inst_621.INIT_2 = 16'h0000;
defparam ram16sdp_inst_621.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_622 (
    .DO(ram16sdp_inst_622_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_233),
    .CLK(clk)
);

defparam ram16sdp_inst_622.INIT_0 = 16'h0000;
defparam ram16sdp_inst_622.INIT_1 = 16'h0000;
defparam ram16sdp_inst_622.INIT_2 = 16'h0000;
defparam ram16sdp_inst_622.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_623 (
    .DO(ram16sdp_inst_623_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_233),
    .CLK(clk)
);

defparam ram16sdp_inst_623.INIT_0 = 16'h0000;
defparam ram16sdp_inst_623.INIT_1 = 16'h0000;
defparam ram16sdp_inst_623.INIT_2 = 16'h0000;
defparam ram16sdp_inst_623.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_624 (
    .DO(ram16sdp_inst_624_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_236),
    .CLK(clk)
);

defparam ram16sdp_inst_624.INIT_0 = 16'h0000;
defparam ram16sdp_inst_624.INIT_1 = 16'h0000;
defparam ram16sdp_inst_624.INIT_2 = 16'h0000;
defparam ram16sdp_inst_624.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_625 (
    .DO(ram16sdp_inst_625_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_236),
    .CLK(clk)
);

defparam ram16sdp_inst_625.INIT_0 = 16'h0000;
defparam ram16sdp_inst_625.INIT_1 = 16'h0000;
defparam ram16sdp_inst_625.INIT_2 = 16'h0000;
defparam ram16sdp_inst_625.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_626 (
    .DO(ram16sdp_inst_626_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_236),
    .CLK(clk)
);

defparam ram16sdp_inst_626.INIT_0 = 16'h0000;
defparam ram16sdp_inst_626.INIT_1 = 16'h0000;
defparam ram16sdp_inst_626.INIT_2 = 16'h0000;
defparam ram16sdp_inst_626.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_627 (
    .DO(ram16sdp_inst_627_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_236),
    .CLK(clk)
);

defparam ram16sdp_inst_627.INIT_0 = 16'h0000;
defparam ram16sdp_inst_627.INIT_1 = 16'h0000;
defparam ram16sdp_inst_627.INIT_2 = 16'h0000;
defparam ram16sdp_inst_627.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_628 (
    .DO(ram16sdp_inst_628_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_236),
    .CLK(clk)
);

defparam ram16sdp_inst_628.INIT_0 = 16'h0000;
defparam ram16sdp_inst_628.INIT_1 = 16'h0000;
defparam ram16sdp_inst_628.INIT_2 = 16'h0000;
defparam ram16sdp_inst_628.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_629 (
    .DO(ram16sdp_inst_629_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_236),
    .CLK(clk)
);

defparam ram16sdp_inst_629.INIT_0 = 16'h0000;
defparam ram16sdp_inst_629.INIT_1 = 16'h0000;
defparam ram16sdp_inst_629.INIT_2 = 16'h0000;
defparam ram16sdp_inst_629.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_630 (
    .DO(ram16sdp_inst_630_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_236),
    .CLK(clk)
);

defparam ram16sdp_inst_630.INIT_0 = 16'h0000;
defparam ram16sdp_inst_630.INIT_1 = 16'h0000;
defparam ram16sdp_inst_630.INIT_2 = 16'h0000;
defparam ram16sdp_inst_630.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_631 (
    .DO(ram16sdp_inst_631_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_236),
    .CLK(clk)
);

defparam ram16sdp_inst_631.INIT_0 = 16'h0000;
defparam ram16sdp_inst_631.INIT_1 = 16'h0000;
defparam ram16sdp_inst_631.INIT_2 = 16'h0000;
defparam ram16sdp_inst_631.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_632 (
    .DO(ram16sdp_inst_632_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16sdp_inst_632.INIT_0 = 16'h0000;
defparam ram16sdp_inst_632.INIT_1 = 16'h0000;
defparam ram16sdp_inst_632.INIT_2 = 16'h0000;
defparam ram16sdp_inst_632.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_633 (
    .DO(ram16sdp_inst_633_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16sdp_inst_633.INIT_0 = 16'h0000;
defparam ram16sdp_inst_633.INIT_1 = 16'h0000;
defparam ram16sdp_inst_633.INIT_2 = 16'h0000;
defparam ram16sdp_inst_633.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_634 (
    .DO(ram16sdp_inst_634_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16sdp_inst_634.INIT_0 = 16'h0000;
defparam ram16sdp_inst_634.INIT_1 = 16'h0000;
defparam ram16sdp_inst_634.INIT_2 = 16'h0000;
defparam ram16sdp_inst_634.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_635 (
    .DO(ram16sdp_inst_635_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16sdp_inst_635.INIT_0 = 16'h0000;
defparam ram16sdp_inst_635.INIT_1 = 16'h0000;
defparam ram16sdp_inst_635.INIT_2 = 16'h0000;
defparam ram16sdp_inst_635.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_636 (
    .DO(ram16sdp_inst_636_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16sdp_inst_636.INIT_0 = 16'h0000;
defparam ram16sdp_inst_636.INIT_1 = 16'h0000;
defparam ram16sdp_inst_636.INIT_2 = 16'h0000;
defparam ram16sdp_inst_636.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_637 (
    .DO(ram16sdp_inst_637_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16sdp_inst_637.INIT_0 = 16'h0000;
defparam ram16sdp_inst_637.INIT_1 = 16'h0000;
defparam ram16sdp_inst_637.INIT_2 = 16'h0000;
defparam ram16sdp_inst_637.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_638 (
    .DO(ram16sdp_inst_638_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16sdp_inst_638.INIT_0 = 16'h0000;
defparam ram16sdp_inst_638.INIT_1 = 16'h0000;
defparam ram16sdp_inst_638.INIT_2 = 16'h0000;
defparam ram16sdp_inst_638.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_639 (
    .DO(ram16sdp_inst_639_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16sdp_inst_639.INIT_0 = 16'h0000;
defparam ram16sdp_inst_639.INIT_1 = 16'h0000;
defparam ram16sdp_inst_639.INIT_2 = 16'h0000;
defparam ram16sdp_inst_639.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_640 (
    .DO(ram16sdp_inst_640_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_242),
    .CLK(clk)
);

defparam ram16sdp_inst_640.INIT_0 = 16'h0000;
defparam ram16sdp_inst_640.INIT_1 = 16'h0000;
defparam ram16sdp_inst_640.INIT_2 = 16'h0000;
defparam ram16sdp_inst_640.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_641 (
    .DO(ram16sdp_inst_641_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_242),
    .CLK(clk)
);

defparam ram16sdp_inst_641.INIT_0 = 16'h0000;
defparam ram16sdp_inst_641.INIT_1 = 16'h0000;
defparam ram16sdp_inst_641.INIT_2 = 16'h0000;
defparam ram16sdp_inst_641.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_642 (
    .DO(ram16sdp_inst_642_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_242),
    .CLK(clk)
);

defparam ram16sdp_inst_642.INIT_0 = 16'h0000;
defparam ram16sdp_inst_642.INIT_1 = 16'h0000;
defparam ram16sdp_inst_642.INIT_2 = 16'h0000;
defparam ram16sdp_inst_642.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_643 (
    .DO(ram16sdp_inst_643_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_242),
    .CLK(clk)
);

defparam ram16sdp_inst_643.INIT_0 = 16'h0000;
defparam ram16sdp_inst_643.INIT_1 = 16'h0000;
defparam ram16sdp_inst_643.INIT_2 = 16'h0000;
defparam ram16sdp_inst_643.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_644 (
    .DO(ram16sdp_inst_644_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_242),
    .CLK(clk)
);

defparam ram16sdp_inst_644.INIT_0 = 16'h0000;
defparam ram16sdp_inst_644.INIT_1 = 16'h0000;
defparam ram16sdp_inst_644.INIT_2 = 16'h0000;
defparam ram16sdp_inst_644.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_645 (
    .DO(ram16sdp_inst_645_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_242),
    .CLK(clk)
);

defparam ram16sdp_inst_645.INIT_0 = 16'h0000;
defparam ram16sdp_inst_645.INIT_1 = 16'h0000;
defparam ram16sdp_inst_645.INIT_2 = 16'h0000;
defparam ram16sdp_inst_645.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_646 (
    .DO(ram16sdp_inst_646_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_242),
    .CLK(clk)
);

defparam ram16sdp_inst_646.INIT_0 = 16'h0000;
defparam ram16sdp_inst_646.INIT_1 = 16'h0000;
defparam ram16sdp_inst_646.INIT_2 = 16'h0000;
defparam ram16sdp_inst_646.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_647 (
    .DO(ram16sdp_inst_647_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_242),
    .CLK(clk)
);

defparam ram16sdp_inst_647.INIT_0 = 16'h0000;
defparam ram16sdp_inst_647.INIT_1 = 16'h0000;
defparam ram16sdp_inst_647.INIT_2 = 16'h0000;
defparam ram16sdp_inst_647.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_648 (
    .DO(ram16sdp_inst_648_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_245),
    .CLK(clk)
);

defparam ram16sdp_inst_648.INIT_0 = 16'h0000;
defparam ram16sdp_inst_648.INIT_1 = 16'h0000;
defparam ram16sdp_inst_648.INIT_2 = 16'h0000;
defparam ram16sdp_inst_648.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_649 (
    .DO(ram16sdp_inst_649_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_245),
    .CLK(clk)
);

defparam ram16sdp_inst_649.INIT_0 = 16'h0000;
defparam ram16sdp_inst_649.INIT_1 = 16'h0000;
defparam ram16sdp_inst_649.INIT_2 = 16'h0000;
defparam ram16sdp_inst_649.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_650 (
    .DO(ram16sdp_inst_650_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_245),
    .CLK(clk)
);

defparam ram16sdp_inst_650.INIT_0 = 16'h0000;
defparam ram16sdp_inst_650.INIT_1 = 16'h0000;
defparam ram16sdp_inst_650.INIT_2 = 16'h0000;
defparam ram16sdp_inst_650.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_651 (
    .DO(ram16sdp_inst_651_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_245),
    .CLK(clk)
);

defparam ram16sdp_inst_651.INIT_0 = 16'h0000;
defparam ram16sdp_inst_651.INIT_1 = 16'h0000;
defparam ram16sdp_inst_651.INIT_2 = 16'h0000;
defparam ram16sdp_inst_651.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_652 (
    .DO(ram16sdp_inst_652_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_245),
    .CLK(clk)
);

defparam ram16sdp_inst_652.INIT_0 = 16'h0000;
defparam ram16sdp_inst_652.INIT_1 = 16'h0000;
defparam ram16sdp_inst_652.INIT_2 = 16'h0000;
defparam ram16sdp_inst_652.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_653 (
    .DO(ram16sdp_inst_653_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_245),
    .CLK(clk)
);

defparam ram16sdp_inst_653.INIT_0 = 16'h0000;
defparam ram16sdp_inst_653.INIT_1 = 16'h0000;
defparam ram16sdp_inst_653.INIT_2 = 16'h0000;
defparam ram16sdp_inst_653.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_654 (
    .DO(ram16sdp_inst_654_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_245),
    .CLK(clk)
);

defparam ram16sdp_inst_654.INIT_0 = 16'h0000;
defparam ram16sdp_inst_654.INIT_1 = 16'h0000;
defparam ram16sdp_inst_654.INIT_2 = 16'h0000;
defparam ram16sdp_inst_654.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_655 (
    .DO(ram16sdp_inst_655_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_245),
    .CLK(clk)
);

defparam ram16sdp_inst_655.INIT_0 = 16'h0000;
defparam ram16sdp_inst_655.INIT_1 = 16'h0000;
defparam ram16sdp_inst_655.INIT_2 = 16'h0000;
defparam ram16sdp_inst_655.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_656 (
    .DO(ram16sdp_inst_656_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_248),
    .CLK(clk)
);

defparam ram16sdp_inst_656.INIT_0 = 16'h0000;
defparam ram16sdp_inst_656.INIT_1 = 16'h0000;
defparam ram16sdp_inst_656.INIT_2 = 16'h0000;
defparam ram16sdp_inst_656.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_657 (
    .DO(ram16sdp_inst_657_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_248),
    .CLK(clk)
);

defparam ram16sdp_inst_657.INIT_0 = 16'h0000;
defparam ram16sdp_inst_657.INIT_1 = 16'h0000;
defparam ram16sdp_inst_657.INIT_2 = 16'h0000;
defparam ram16sdp_inst_657.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_658 (
    .DO(ram16sdp_inst_658_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_248),
    .CLK(clk)
);

defparam ram16sdp_inst_658.INIT_0 = 16'h0000;
defparam ram16sdp_inst_658.INIT_1 = 16'h0000;
defparam ram16sdp_inst_658.INIT_2 = 16'h0000;
defparam ram16sdp_inst_658.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_659 (
    .DO(ram16sdp_inst_659_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_248),
    .CLK(clk)
);

defparam ram16sdp_inst_659.INIT_0 = 16'h0000;
defparam ram16sdp_inst_659.INIT_1 = 16'h0000;
defparam ram16sdp_inst_659.INIT_2 = 16'h0000;
defparam ram16sdp_inst_659.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_660 (
    .DO(ram16sdp_inst_660_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_248),
    .CLK(clk)
);

defparam ram16sdp_inst_660.INIT_0 = 16'h0000;
defparam ram16sdp_inst_660.INIT_1 = 16'h0000;
defparam ram16sdp_inst_660.INIT_2 = 16'h0000;
defparam ram16sdp_inst_660.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_661 (
    .DO(ram16sdp_inst_661_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_248),
    .CLK(clk)
);

defparam ram16sdp_inst_661.INIT_0 = 16'h0000;
defparam ram16sdp_inst_661.INIT_1 = 16'h0000;
defparam ram16sdp_inst_661.INIT_2 = 16'h0000;
defparam ram16sdp_inst_661.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_662 (
    .DO(ram16sdp_inst_662_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_248),
    .CLK(clk)
);

defparam ram16sdp_inst_662.INIT_0 = 16'h0000;
defparam ram16sdp_inst_662.INIT_1 = 16'h0000;
defparam ram16sdp_inst_662.INIT_2 = 16'h0000;
defparam ram16sdp_inst_662.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_663 (
    .DO(ram16sdp_inst_663_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_248),
    .CLK(clk)
);

defparam ram16sdp_inst_663.INIT_0 = 16'h0000;
defparam ram16sdp_inst_663.INIT_1 = 16'h0000;
defparam ram16sdp_inst_663.INIT_2 = 16'h0000;
defparam ram16sdp_inst_663.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_664 (
    .DO(ram16sdp_inst_664_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16sdp_inst_664.INIT_0 = 16'h0000;
defparam ram16sdp_inst_664.INIT_1 = 16'h0000;
defparam ram16sdp_inst_664.INIT_2 = 16'h0000;
defparam ram16sdp_inst_664.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_665 (
    .DO(ram16sdp_inst_665_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16sdp_inst_665.INIT_0 = 16'h0000;
defparam ram16sdp_inst_665.INIT_1 = 16'h0000;
defparam ram16sdp_inst_665.INIT_2 = 16'h0000;
defparam ram16sdp_inst_665.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_666 (
    .DO(ram16sdp_inst_666_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16sdp_inst_666.INIT_0 = 16'h0000;
defparam ram16sdp_inst_666.INIT_1 = 16'h0000;
defparam ram16sdp_inst_666.INIT_2 = 16'h0000;
defparam ram16sdp_inst_666.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_667 (
    .DO(ram16sdp_inst_667_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16sdp_inst_667.INIT_0 = 16'h0000;
defparam ram16sdp_inst_667.INIT_1 = 16'h0000;
defparam ram16sdp_inst_667.INIT_2 = 16'h0000;
defparam ram16sdp_inst_667.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_668 (
    .DO(ram16sdp_inst_668_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16sdp_inst_668.INIT_0 = 16'h0000;
defparam ram16sdp_inst_668.INIT_1 = 16'h0000;
defparam ram16sdp_inst_668.INIT_2 = 16'h0000;
defparam ram16sdp_inst_668.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_669 (
    .DO(ram16sdp_inst_669_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16sdp_inst_669.INIT_0 = 16'h0000;
defparam ram16sdp_inst_669.INIT_1 = 16'h0000;
defparam ram16sdp_inst_669.INIT_2 = 16'h0000;
defparam ram16sdp_inst_669.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_670 (
    .DO(ram16sdp_inst_670_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16sdp_inst_670.INIT_0 = 16'h0000;
defparam ram16sdp_inst_670.INIT_1 = 16'h0000;
defparam ram16sdp_inst_670.INIT_2 = 16'h0000;
defparam ram16sdp_inst_670.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_671 (
    .DO(ram16sdp_inst_671_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16sdp_inst_671.INIT_0 = 16'h0000;
defparam ram16sdp_inst_671.INIT_1 = 16'h0000;
defparam ram16sdp_inst_671.INIT_2 = 16'h0000;
defparam ram16sdp_inst_671.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_672 (
    .DO(ram16sdp_inst_672_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_254),
    .CLK(clk)
);

defparam ram16sdp_inst_672.INIT_0 = 16'h0000;
defparam ram16sdp_inst_672.INIT_1 = 16'h0000;
defparam ram16sdp_inst_672.INIT_2 = 16'h0000;
defparam ram16sdp_inst_672.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_673 (
    .DO(ram16sdp_inst_673_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_254),
    .CLK(clk)
);

defparam ram16sdp_inst_673.INIT_0 = 16'h0000;
defparam ram16sdp_inst_673.INIT_1 = 16'h0000;
defparam ram16sdp_inst_673.INIT_2 = 16'h0000;
defparam ram16sdp_inst_673.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_674 (
    .DO(ram16sdp_inst_674_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_254),
    .CLK(clk)
);

defparam ram16sdp_inst_674.INIT_0 = 16'h0000;
defparam ram16sdp_inst_674.INIT_1 = 16'h0000;
defparam ram16sdp_inst_674.INIT_2 = 16'h0000;
defparam ram16sdp_inst_674.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_675 (
    .DO(ram16sdp_inst_675_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_254),
    .CLK(clk)
);

defparam ram16sdp_inst_675.INIT_0 = 16'h0000;
defparam ram16sdp_inst_675.INIT_1 = 16'h0000;
defparam ram16sdp_inst_675.INIT_2 = 16'h0000;
defparam ram16sdp_inst_675.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_676 (
    .DO(ram16sdp_inst_676_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_254),
    .CLK(clk)
);

defparam ram16sdp_inst_676.INIT_0 = 16'h0000;
defparam ram16sdp_inst_676.INIT_1 = 16'h0000;
defparam ram16sdp_inst_676.INIT_2 = 16'h0000;
defparam ram16sdp_inst_676.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_677 (
    .DO(ram16sdp_inst_677_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_254),
    .CLK(clk)
);

defparam ram16sdp_inst_677.INIT_0 = 16'h0000;
defparam ram16sdp_inst_677.INIT_1 = 16'h0000;
defparam ram16sdp_inst_677.INIT_2 = 16'h0000;
defparam ram16sdp_inst_677.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_678 (
    .DO(ram16sdp_inst_678_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_254),
    .CLK(clk)
);

defparam ram16sdp_inst_678.INIT_0 = 16'h0000;
defparam ram16sdp_inst_678.INIT_1 = 16'h0000;
defparam ram16sdp_inst_678.INIT_2 = 16'h0000;
defparam ram16sdp_inst_678.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_679 (
    .DO(ram16sdp_inst_679_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_254),
    .CLK(clk)
);

defparam ram16sdp_inst_679.INIT_0 = 16'h0000;
defparam ram16sdp_inst_679.INIT_1 = 16'h0000;
defparam ram16sdp_inst_679.INIT_2 = 16'h0000;
defparam ram16sdp_inst_679.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_680 (
    .DO(ram16sdp_inst_680_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_257),
    .CLK(clk)
);

defparam ram16sdp_inst_680.INIT_0 = 16'h0000;
defparam ram16sdp_inst_680.INIT_1 = 16'h0000;
defparam ram16sdp_inst_680.INIT_2 = 16'h0000;
defparam ram16sdp_inst_680.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_681 (
    .DO(ram16sdp_inst_681_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_257),
    .CLK(clk)
);

defparam ram16sdp_inst_681.INIT_0 = 16'h0000;
defparam ram16sdp_inst_681.INIT_1 = 16'h0000;
defparam ram16sdp_inst_681.INIT_2 = 16'h0000;
defparam ram16sdp_inst_681.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_682 (
    .DO(ram16sdp_inst_682_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_257),
    .CLK(clk)
);

defparam ram16sdp_inst_682.INIT_0 = 16'h0000;
defparam ram16sdp_inst_682.INIT_1 = 16'h0000;
defparam ram16sdp_inst_682.INIT_2 = 16'h0000;
defparam ram16sdp_inst_682.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_683 (
    .DO(ram16sdp_inst_683_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_257),
    .CLK(clk)
);

defparam ram16sdp_inst_683.INIT_0 = 16'h0000;
defparam ram16sdp_inst_683.INIT_1 = 16'h0000;
defparam ram16sdp_inst_683.INIT_2 = 16'h0000;
defparam ram16sdp_inst_683.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_684 (
    .DO(ram16sdp_inst_684_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_257),
    .CLK(clk)
);

defparam ram16sdp_inst_684.INIT_0 = 16'h0000;
defparam ram16sdp_inst_684.INIT_1 = 16'h0000;
defparam ram16sdp_inst_684.INIT_2 = 16'h0000;
defparam ram16sdp_inst_684.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_685 (
    .DO(ram16sdp_inst_685_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_257),
    .CLK(clk)
);

defparam ram16sdp_inst_685.INIT_0 = 16'h0000;
defparam ram16sdp_inst_685.INIT_1 = 16'h0000;
defparam ram16sdp_inst_685.INIT_2 = 16'h0000;
defparam ram16sdp_inst_685.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_686 (
    .DO(ram16sdp_inst_686_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_257),
    .CLK(clk)
);

defparam ram16sdp_inst_686.INIT_0 = 16'h0000;
defparam ram16sdp_inst_686.INIT_1 = 16'h0000;
defparam ram16sdp_inst_686.INIT_2 = 16'h0000;
defparam ram16sdp_inst_686.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_687 (
    .DO(ram16sdp_inst_687_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_257),
    .CLK(clk)
);

defparam ram16sdp_inst_687.INIT_0 = 16'h0000;
defparam ram16sdp_inst_687.INIT_1 = 16'h0000;
defparam ram16sdp_inst_687.INIT_2 = 16'h0000;
defparam ram16sdp_inst_687.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_688 (
    .DO(ram16sdp_inst_688_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_260),
    .CLK(clk)
);

defparam ram16sdp_inst_688.INIT_0 = 16'h0000;
defparam ram16sdp_inst_688.INIT_1 = 16'h0000;
defparam ram16sdp_inst_688.INIT_2 = 16'h0000;
defparam ram16sdp_inst_688.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_689 (
    .DO(ram16sdp_inst_689_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_260),
    .CLK(clk)
);

defparam ram16sdp_inst_689.INIT_0 = 16'h0000;
defparam ram16sdp_inst_689.INIT_1 = 16'h0000;
defparam ram16sdp_inst_689.INIT_2 = 16'h0000;
defparam ram16sdp_inst_689.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_690 (
    .DO(ram16sdp_inst_690_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_260),
    .CLK(clk)
);

defparam ram16sdp_inst_690.INIT_0 = 16'h0000;
defparam ram16sdp_inst_690.INIT_1 = 16'h0000;
defparam ram16sdp_inst_690.INIT_2 = 16'h0000;
defparam ram16sdp_inst_690.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_691 (
    .DO(ram16sdp_inst_691_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_260),
    .CLK(clk)
);

defparam ram16sdp_inst_691.INIT_0 = 16'h0000;
defparam ram16sdp_inst_691.INIT_1 = 16'h0000;
defparam ram16sdp_inst_691.INIT_2 = 16'h0000;
defparam ram16sdp_inst_691.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_692 (
    .DO(ram16sdp_inst_692_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_260),
    .CLK(clk)
);

defparam ram16sdp_inst_692.INIT_0 = 16'h0000;
defparam ram16sdp_inst_692.INIT_1 = 16'h0000;
defparam ram16sdp_inst_692.INIT_2 = 16'h0000;
defparam ram16sdp_inst_692.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_693 (
    .DO(ram16sdp_inst_693_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_260),
    .CLK(clk)
);

defparam ram16sdp_inst_693.INIT_0 = 16'h0000;
defparam ram16sdp_inst_693.INIT_1 = 16'h0000;
defparam ram16sdp_inst_693.INIT_2 = 16'h0000;
defparam ram16sdp_inst_693.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_694 (
    .DO(ram16sdp_inst_694_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_260),
    .CLK(clk)
);

defparam ram16sdp_inst_694.INIT_0 = 16'h0000;
defparam ram16sdp_inst_694.INIT_1 = 16'h0000;
defparam ram16sdp_inst_694.INIT_2 = 16'h0000;
defparam ram16sdp_inst_694.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_695 (
    .DO(ram16sdp_inst_695_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_260),
    .CLK(clk)
);

defparam ram16sdp_inst_695.INIT_0 = 16'h0000;
defparam ram16sdp_inst_695.INIT_1 = 16'h0000;
defparam ram16sdp_inst_695.INIT_2 = 16'h0000;
defparam ram16sdp_inst_695.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_696 (
    .DO(ram16sdp_inst_696_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16sdp_inst_696.INIT_0 = 16'h0000;
defparam ram16sdp_inst_696.INIT_1 = 16'h0000;
defparam ram16sdp_inst_696.INIT_2 = 16'h0000;
defparam ram16sdp_inst_696.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_697 (
    .DO(ram16sdp_inst_697_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16sdp_inst_697.INIT_0 = 16'h0000;
defparam ram16sdp_inst_697.INIT_1 = 16'h0000;
defparam ram16sdp_inst_697.INIT_2 = 16'h0000;
defparam ram16sdp_inst_697.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_698 (
    .DO(ram16sdp_inst_698_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16sdp_inst_698.INIT_0 = 16'h0000;
defparam ram16sdp_inst_698.INIT_1 = 16'h0000;
defparam ram16sdp_inst_698.INIT_2 = 16'h0000;
defparam ram16sdp_inst_698.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_699 (
    .DO(ram16sdp_inst_699_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16sdp_inst_699.INIT_0 = 16'h0000;
defparam ram16sdp_inst_699.INIT_1 = 16'h0000;
defparam ram16sdp_inst_699.INIT_2 = 16'h0000;
defparam ram16sdp_inst_699.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_700 (
    .DO(ram16sdp_inst_700_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16sdp_inst_700.INIT_0 = 16'h0000;
defparam ram16sdp_inst_700.INIT_1 = 16'h0000;
defparam ram16sdp_inst_700.INIT_2 = 16'h0000;
defparam ram16sdp_inst_700.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_701 (
    .DO(ram16sdp_inst_701_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16sdp_inst_701.INIT_0 = 16'h0000;
defparam ram16sdp_inst_701.INIT_1 = 16'h0000;
defparam ram16sdp_inst_701.INIT_2 = 16'h0000;
defparam ram16sdp_inst_701.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_702 (
    .DO(ram16sdp_inst_702_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16sdp_inst_702.INIT_0 = 16'h0000;
defparam ram16sdp_inst_702.INIT_1 = 16'h0000;
defparam ram16sdp_inst_702.INIT_2 = 16'h0000;
defparam ram16sdp_inst_702.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_703 (
    .DO(ram16sdp_inst_703_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16sdp_inst_703.INIT_0 = 16'h0000;
defparam ram16sdp_inst_703.INIT_1 = 16'h0000;
defparam ram16sdp_inst_703.INIT_2 = 16'h0000;
defparam ram16sdp_inst_703.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_704 (
    .DO(ram16sdp_inst_704_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_266),
    .CLK(clk)
);

defparam ram16sdp_inst_704.INIT_0 = 16'h0000;
defparam ram16sdp_inst_704.INIT_1 = 16'h0000;
defparam ram16sdp_inst_704.INIT_2 = 16'h0000;
defparam ram16sdp_inst_704.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_705 (
    .DO(ram16sdp_inst_705_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_266),
    .CLK(clk)
);

defparam ram16sdp_inst_705.INIT_0 = 16'h0000;
defparam ram16sdp_inst_705.INIT_1 = 16'h0000;
defparam ram16sdp_inst_705.INIT_2 = 16'h0000;
defparam ram16sdp_inst_705.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_706 (
    .DO(ram16sdp_inst_706_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_266),
    .CLK(clk)
);

defparam ram16sdp_inst_706.INIT_0 = 16'h0000;
defparam ram16sdp_inst_706.INIT_1 = 16'h0000;
defparam ram16sdp_inst_706.INIT_2 = 16'h0000;
defparam ram16sdp_inst_706.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_707 (
    .DO(ram16sdp_inst_707_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_266),
    .CLK(clk)
);

defparam ram16sdp_inst_707.INIT_0 = 16'h0000;
defparam ram16sdp_inst_707.INIT_1 = 16'h0000;
defparam ram16sdp_inst_707.INIT_2 = 16'h0000;
defparam ram16sdp_inst_707.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_708 (
    .DO(ram16sdp_inst_708_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_266),
    .CLK(clk)
);

defparam ram16sdp_inst_708.INIT_0 = 16'h0000;
defparam ram16sdp_inst_708.INIT_1 = 16'h0000;
defparam ram16sdp_inst_708.INIT_2 = 16'h0000;
defparam ram16sdp_inst_708.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_709 (
    .DO(ram16sdp_inst_709_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_266),
    .CLK(clk)
);

defparam ram16sdp_inst_709.INIT_0 = 16'h0000;
defparam ram16sdp_inst_709.INIT_1 = 16'h0000;
defparam ram16sdp_inst_709.INIT_2 = 16'h0000;
defparam ram16sdp_inst_709.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_710 (
    .DO(ram16sdp_inst_710_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_266),
    .CLK(clk)
);

defparam ram16sdp_inst_710.INIT_0 = 16'h0000;
defparam ram16sdp_inst_710.INIT_1 = 16'h0000;
defparam ram16sdp_inst_710.INIT_2 = 16'h0000;
defparam ram16sdp_inst_710.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_711 (
    .DO(ram16sdp_inst_711_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_266),
    .CLK(clk)
);

defparam ram16sdp_inst_711.INIT_0 = 16'h0000;
defparam ram16sdp_inst_711.INIT_1 = 16'h0000;
defparam ram16sdp_inst_711.INIT_2 = 16'h0000;
defparam ram16sdp_inst_711.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_712 (
    .DO(ram16sdp_inst_712_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_269),
    .CLK(clk)
);

defparam ram16sdp_inst_712.INIT_0 = 16'h0000;
defparam ram16sdp_inst_712.INIT_1 = 16'h0000;
defparam ram16sdp_inst_712.INIT_2 = 16'h0000;
defparam ram16sdp_inst_712.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_713 (
    .DO(ram16sdp_inst_713_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_269),
    .CLK(clk)
);

defparam ram16sdp_inst_713.INIT_0 = 16'h0000;
defparam ram16sdp_inst_713.INIT_1 = 16'h0000;
defparam ram16sdp_inst_713.INIT_2 = 16'h0000;
defparam ram16sdp_inst_713.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_714 (
    .DO(ram16sdp_inst_714_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_269),
    .CLK(clk)
);

defparam ram16sdp_inst_714.INIT_0 = 16'h0000;
defparam ram16sdp_inst_714.INIT_1 = 16'h0000;
defparam ram16sdp_inst_714.INIT_2 = 16'h0000;
defparam ram16sdp_inst_714.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_715 (
    .DO(ram16sdp_inst_715_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_269),
    .CLK(clk)
);

defparam ram16sdp_inst_715.INIT_0 = 16'h0000;
defparam ram16sdp_inst_715.INIT_1 = 16'h0000;
defparam ram16sdp_inst_715.INIT_2 = 16'h0000;
defparam ram16sdp_inst_715.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_716 (
    .DO(ram16sdp_inst_716_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_269),
    .CLK(clk)
);

defparam ram16sdp_inst_716.INIT_0 = 16'h0000;
defparam ram16sdp_inst_716.INIT_1 = 16'h0000;
defparam ram16sdp_inst_716.INIT_2 = 16'h0000;
defparam ram16sdp_inst_716.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_717 (
    .DO(ram16sdp_inst_717_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_269),
    .CLK(clk)
);

defparam ram16sdp_inst_717.INIT_0 = 16'h0000;
defparam ram16sdp_inst_717.INIT_1 = 16'h0000;
defparam ram16sdp_inst_717.INIT_2 = 16'h0000;
defparam ram16sdp_inst_717.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_718 (
    .DO(ram16sdp_inst_718_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_269),
    .CLK(clk)
);

defparam ram16sdp_inst_718.INIT_0 = 16'h0000;
defparam ram16sdp_inst_718.INIT_1 = 16'h0000;
defparam ram16sdp_inst_718.INIT_2 = 16'h0000;
defparam ram16sdp_inst_718.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_719 (
    .DO(ram16sdp_inst_719_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_269),
    .CLK(clk)
);

defparam ram16sdp_inst_719.INIT_0 = 16'h0000;
defparam ram16sdp_inst_719.INIT_1 = 16'h0000;
defparam ram16sdp_inst_719.INIT_2 = 16'h0000;
defparam ram16sdp_inst_719.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_720 (
    .DO(ram16sdp_inst_720_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_272),
    .CLK(clk)
);

defparam ram16sdp_inst_720.INIT_0 = 16'h0000;
defparam ram16sdp_inst_720.INIT_1 = 16'h0000;
defparam ram16sdp_inst_720.INIT_2 = 16'h0000;
defparam ram16sdp_inst_720.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_721 (
    .DO(ram16sdp_inst_721_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_272),
    .CLK(clk)
);

defparam ram16sdp_inst_721.INIT_0 = 16'h0000;
defparam ram16sdp_inst_721.INIT_1 = 16'h0000;
defparam ram16sdp_inst_721.INIT_2 = 16'h0000;
defparam ram16sdp_inst_721.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_722 (
    .DO(ram16sdp_inst_722_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_272),
    .CLK(clk)
);

defparam ram16sdp_inst_722.INIT_0 = 16'h0000;
defparam ram16sdp_inst_722.INIT_1 = 16'h0000;
defparam ram16sdp_inst_722.INIT_2 = 16'h0000;
defparam ram16sdp_inst_722.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_723 (
    .DO(ram16sdp_inst_723_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_272),
    .CLK(clk)
);

defparam ram16sdp_inst_723.INIT_0 = 16'h0000;
defparam ram16sdp_inst_723.INIT_1 = 16'h0000;
defparam ram16sdp_inst_723.INIT_2 = 16'h0000;
defparam ram16sdp_inst_723.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_724 (
    .DO(ram16sdp_inst_724_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_272),
    .CLK(clk)
);

defparam ram16sdp_inst_724.INIT_0 = 16'h0000;
defparam ram16sdp_inst_724.INIT_1 = 16'h0000;
defparam ram16sdp_inst_724.INIT_2 = 16'h0000;
defparam ram16sdp_inst_724.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_725 (
    .DO(ram16sdp_inst_725_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_272),
    .CLK(clk)
);

defparam ram16sdp_inst_725.INIT_0 = 16'h0000;
defparam ram16sdp_inst_725.INIT_1 = 16'h0000;
defparam ram16sdp_inst_725.INIT_2 = 16'h0000;
defparam ram16sdp_inst_725.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_726 (
    .DO(ram16sdp_inst_726_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_272),
    .CLK(clk)
);

defparam ram16sdp_inst_726.INIT_0 = 16'h0000;
defparam ram16sdp_inst_726.INIT_1 = 16'h0000;
defparam ram16sdp_inst_726.INIT_2 = 16'h0000;
defparam ram16sdp_inst_726.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_727 (
    .DO(ram16sdp_inst_727_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_272),
    .CLK(clk)
);

defparam ram16sdp_inst_727.INIT_0 = 16'h0000;
defparam ram16sdp_inst_727.INIT_1 = 16'h0000;
defparam ram16sdp_inst_727.INIT_2 = 16'h0000;
defparam ram16sdp_inst_727.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_728 (
    .DO(ram16sdp_inst_728_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16sdp_inst_728.INIT_0 = 16'h0000;
defparam ram16sdp_inst_728.INIT_1 = 16'h0000;
defparam ram16sdp_inst_728.INIT_2 = 16'h0000;
defparam ram16sdp_inst_728.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_729 (
    .DO(ram16sdp_inst_729_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16sdp_inst_729.INIT_0 = 16'h0000;
defparam ram16sdp_inst_729.INIT_1 = 16'h0000;
defparam ram16sdp_inst_729.INIT_2 = 16'h0000;
defparam ram16sdp_inst_729.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_730 (
    .DO(ram16sdp_inst_730_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16sdp_inst_730.INIT_0 = 16'h0000;
defparam ram16sdp_inst_730.INIT_1 = 16'h0000;
defparam ram16sdp_inst_730.INIT_2 = 16'h0000;
defparam ram16sdp_inst_730.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_731 (
    .DO(ram16sdp_inst_731_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16sdp_inst_731.INIT_0 = 16'h0000;
defparam ram16sdp_inst_731.INIT_1 = 16'h0000;
defparam ram16sdp_inst_731.INIT_2 = 16'h0000;
defparam ram16sdp_inst_731.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_732 (
    .DO(ram16sdp_inst_732_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16sdp_inst_732.INIT_0 = 16'h0000;
defparam ram16sdp_inst_732.INIT_1 = 16'h0000;
defparam ram16sdp_inst_732.INIT_2 = 16'h0000;
defparam ram16sdp_inst_732.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_733 (
    .DO(ram16sdp_inst_733_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16sdp_inst_733.INIT_0 = 16'h0000;
defparam ram16sdp_inst_733.INIT_1 = 16'h0000;
defparam ram16sdp_inst_733.INIT_2 = 16'h0000;
defparam ram16sdp_inst_733.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_734 (
    .DO(ram16sdp_inst_734_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16sdp_inst_734.INIT_0 = 16'h0000;
defparam ram16sdp_inst_734.INIT_1 = 16'h0000;
defparam ram16sdp_inst_734.INIT_2 = 16'h0000;
defparam ram16sdp_inst_734.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_735 (
    .DO(ram16sdp_inst_735_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16sdp_inst_735.INIT_0 = 16'h0000;
defparam ram16sdp_inst_735.INIT_1 = 16'h0000;
defparam ram16sdp_inst_735.INIT_2 = 16'h0000;
defparam ram16sdp_inst_735.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_736 (
    .DO(ram16sdp_inst_736_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_278),
    .CLK(clk)
);

defparam ram16sdp_inst_736.INIT_0 = 16'h0000;
defparam ram16sdp_inst_736.INIT_1 = 16'h0000;
defparam ram16sdp_inst_736.INIT_2 = 16'h0000;
defparam ram16sdp_inst_736.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_737 (
    .DO(ram16sdp_inst_737_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_278),
    .CLK(clk)
);

defparam ram16sdp_inst_737.INIT_0 = 16'h0000;
defparam ram16sdp_inst_737.INIT_1 = 16'h0000;
defparam ram16sdp_inst_737.INIT_2 = 16'h0000;
defparam ram16sdp_inst_737.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_738 (
    .DO(ram16sdp_inst_738_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_278),
    .CLK(clk)
);

defparam ram16sdp_inst_738.INIT_0 = 16'h0000;
defparam ram16sdp_inst_738.INIT_1 = 16'h0000;
defparam ram16sdp_inst_738.INIT_2 = 16'h0000;
defparam ram16sdp_inst_738.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_739 (
    .DO(ram16sdp_inst_739_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_278),
    .CLK(clk)
);

defparam ram16sdp_inst_739.INIT_0 = 16'h0000;
defparam ram16sdp_inst_739.INIT_1 = 16'h0000;
defparam ram16sdp_inst_739.INIT_2 = 16'h0000;
defparam ram16sdp_inst_739.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_740 (
    .DO(ram16sdp_inst_740_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_278),
    .CLK(clk)
);

defparam ram16sdp_inst_740.INIT_0 = 16'h0000;
defparam ram16sdp_inst_740.INIT_1 = 16'h0000;
defparam ram16sdp_inst_740.INIT_2 = 16'h0000;
defparam ram16sdp_inst_740.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_741 (
    .DO(ram16sdp_inst_741_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_278),
    .CLK(clk)
);

defparam ram16sdp_inst_741.INIT_0 = 16'h0000;
defparam ram16sdp_inst_741.INIT_1 = 16'h0000;
defparam ram16sdp_inst_741.INIT_2 = 16'h0000;
defparam ram16sdp_inst_741.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_742 (
    .DO(ram16sdp_inst_742_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_278),
    .CLK(clk)
);

defparam ram16sdp_inst_742.INIT_0 = 16'h0000;
defparam ram16sdp_inst_742.INIT_1 = 16'h0000;
defparam ram16sdp_inst_742.INIT_2 = 16'h0000;
defparam ram16sdp_inst_742.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_743 (
    .DO(ram16sdp_inst_743_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_278),
    .CLK(clk)
);

defparam ram16sdp_inst_743.INIT_0 = 16'h0000;
defparam ram16sdp_inst_743.INIT_1 = 16'h0000;
defparam ram16sdp_inst_743.INIT_2 = 16'h0000;
defparam ram16sdp_inst_743.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_744 (
    .DO(ram16sdp_inst_744_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_281),
    .CLK(clk)
);

defparam ram16sdp_inst_744.INIT_0 = 16'h0000;
defparam ram16sdp_inst_744.INIT_1 = 16'h0000;
defparam ram16sdp_inst_744.INIT_2 = 16'h0000;
defparam ram16sdp_inst_744.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_745 (
    .DO(ram16sdp_inst_745_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_281),
    .CLK(clk)
);

defparam ram16sdp_inst_745.INIT_0 = 16'h0000;
defparam ram16sdp_inst_745.INIT_1 = 16'h0000;
defparam ram16sdp_inst_745.INIT_2 = 16'h0000;
defparam ram16sdp_inst_745.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_746 (
    .DO(ram16sdp_inst_746_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_281),
    .CLK(clk)
);

defparam ram16sdp_inst_746.INIT_0 = 16'h0000;
defparam ram16sdp_inst_746.INIT_1 = 16'h0000;
defparam ram16sdp_inst_746.INIT_2 = 16'h0000;
defparam ram16sdp_inst_746.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_747 (
    .DO(ram16sdp_inst_747_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_281),
    .CLK(clk)
);

defparam ram16sdp_inst_747.INIT_0 = 16'h0000;
defparam ram16sdp_inst_747.INIT_1 = 16'h0000;
defparam ram16sdp_inst_747.INIT_2 = 16'h0000;
defparam ram16sdp_inst_747.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_748 (
    .DO(ram16sdp_inst_748_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_281),
    .CLK(clk)
);

defparam ram16sdp_inst_748.INIT_0 = 16'h0000;
defparam ram16sdp_inst_748.INIT_1 = 16'h0000;
defparam ram16sdp_inst_748.INIT_2 = 16'h0000;
defparam ram16sdp_inst_748.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_749 (
    .DO(ram16sdp_inst_749_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_281),
    .CLK(clk)
);

defparam ram16sdp_inst_749.INIT_0 = 16'h0000;
defparam ram16sdp_inst_749.INIT_1 = 16'h0000;
defparam ram16sdp_inst_749.INIT_2 = 16'h0000;
defparam ram16sdp_inst_749.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_750 (
    .DO(ram16sdp_inst_750_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_281),
    .CLK(clk)
);

defparam ram16sdp_inst_750.INIT_0 = 16'h0000;
defparam ram16sdp_inst_750.INIT_1 = 16'h0000;
defparam ram16sdp_inst_750.INIT_2 = 16'h0000;
defparam ram16sdp_inst_750.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_751 (
    .DO(ram16sdp_inst_751_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_281),
    .CLK(clk)
);

defparam ram16sdp_inst_751.INIT_0 = 16'h0000;
defparam ram16sdp_inst_751.INIT_1 = 16'h0000;
defparam ram16sdp_inst_751.INIT_2 = 16'h0000;
defparam ram16sdp_inst_751.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_752 (
    .DO(ram16sdp_inst_752_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_284),
    .CLK(clk)
);

defparam ram16sdp_inst_752.INIT_0 = 16'h0000;
defparam ram16sdp_inst_752.INIT_1 = 16'h0000;
defparam ram16sdp_inst_752.INIT_2 = 16'h0000;
defparam ram16sdp_inst_752.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_753 (
    .DO(ram16sdp_inst_753_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_284),
    .CLK(clk)
);

defparam ram16sdp_inst_753.INIT_0 = 16'h0000;
defparam ram16sdp_inst_753.INIT_1 = 16'h0000;
defparam ram16sdp_inst_753.INIT_2 = 16'h0000;
defparam ram16sdp_inst_753.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_754 (
    .DO(ram16sdp_inst_754_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_284),
    .CLK(clk)
);

defparam ram16sdp_inst_754.INIT_0 = 16'h0000;
defparam ram16sdp_inst_754.INIT_1 = 16'h0000;
defparam ram16sdp_inst_754.INIT_2 = 16'h0000;
defparam ram16sdp_inst_754.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_755 (
    .DO(ram16sdp_inst_755_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_284),
    .CLK(clk)
);

defparam ram16sdp_inst_755.INIT_0 = 16'h0000;
defparam ram16sdp_inst_755.INIT_1 = 16'h0000;
defparam ram16sdp_inst_755.INIT_2 = 16'h0000;
defparam ram16sdp_inst_755.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_756 (
    .DO(ram16sdp_inst_756_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_284),
    .CLK(clk)
);

defparam ram16sdp_inst_756.INIT_0 = 16'h0000;
defparam ram16sdp_inst_756.INIT_1 = 16'h0000;
defparam ram16sdp_inst_756.INIT_2 = 16'h0000;
defparam ram16sdp_inst_756.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_757 (
    .DO(ram16sdp_inst_757_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_284),
    .CLK(clk)
);

defparam ram16sdp_inst_757.INIT_0 = 16'h0000;
defparam ram16sdp_inst_757.INIT_1 = 16'h0000;
defparam ram16sdp_inst_757.INIT_2 = 16'h0000;
defparam ram16sdp_inst_757.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_758 (
    .DO(ram16sdp_inst_758_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_284),
    .CLK(clk)
);

defparam ram16sdp_inst_758.INIT_0 = 16'h0000;
defparam ram16sdp_inst_758.INIT_1 = 16'h0000;
defparam ram16sdp_inst_758.INIT_2 = 16'h0000;
defparam ram16sdp_inst_758.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_759 (
    .DO(ram16sdp_inst_759_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_284),
    .CLK(clk)
);

defparam ram16sdp_inst_759.INIT_0 = 16'h0000;
defparam ram16sdp_inst_759.INIT_1 = 16'h0000;
defparam ram16sdp_inst_759.INIT_2 = 16'h0000;
defparam ram16sdp_inst_759.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_760 (
    .DO(ram16sdp_inst_760_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16sdp_inst_760.INIT_0 = 16'h0000;
defparam ram16sdp_inst_760.INIT_1 = 16'h0000;
defparam ram16sdp_inst_760.INIT_2 = 16'h0000;
defparam ram16sdp_inst_760.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_761 (
    .DO(ram16sdp_inst_761_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16sdp_inst_761.INIT_0 = 16'h0000;
defparam ram16sdp_inst_761.INIT_1 = 16'h0000;
defparam ram16sdp_inst_761.INIT_2 = 16'h0000;
defparam ram16sdp_inst_761.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_762 (
    .DO(ram16sdp_inst_762_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16sdp_inst_762.INIT_0 = 16'h0000;
defparam ram16sdp_inst_762.INIT_1 = 16'h0000;
defparam ram16sdp_inst_762.INIT_2 = 16'h0000;
defparam ram16sdp_inst_762.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_763 (
    .DO(ram16sdp_inst_763_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16sdp_inst_763.INIT_0 = 16'h0000;
defparam ram16sdp_inst_763.INIT_1 = 16'h0000;
defparam ram16sdp_inst_763.INIT_2 = 16'h0000;
defparam ram16sdp_inst_763.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_764 (
    .DO(ram16sdp_inst_764_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16sdp_inst_764.INIT_0 = 16'h0000;
defparam ram16sdp_inst_764.INIT_1 = 16'h0000;
defparam ram16sdp_inst_764.INIT_2 = 16'h0000;
defparam ram16sdp_inst_764.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_765 (
    .DO(ram16sdp_inst_765_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16sdp_inst_765.INIT_0 = 16'h0000;
defparam ram16sdp_inst_765.INIT_1 = 16'h0000;
defparam ram16sdp_inst_765.INIT_2 = 16'h0000;
defparam ram16sdp_inst_765.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_766 (
    .DO(ram16sdp_inst_766_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16sdp_inst_766.INIT_0 = 16'h0000;
defparam ram16sdp_inst_766.INIT_1 = 16'h0000;
defparam ram16sdp_inst_766.INIT_2 = 16'h0000;
defparam ram16sdp_inst_766.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_767 (
    .DO(ram16sdp_inst_767_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16sdp_inst_767.INIT_0 = 16'h0000;
defparam ram16sdp_inst_767.INIT_1 = 16'h0000;
defparam ram16sdp_inst_767.INIT_2 = 16'h0000;
defparam ram16sdp_inst_767.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_768 (
    .DO(ram16sdp_inst_768_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_290),
    .CLK(clk)
);

defparam ram16sdp_inst_768.INIT_0 = 16'h0000;
defparam ram16sdp_inst_768.INIT_1 = 16'h0000;
defparam ram16sdp_inst_768.INIT_2 = 16'h0000;
defparam ram16sdp_inst_768.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_769 (
    .DO(ram16sdp_inst_769_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_290),
    .CLK(clk)
);

defparam ram16sdp_inst_769.INIT_0 = 16'h0000;
defparam ram16sdp_inst_769.INIT_1 = 16'h0000;
defparam ram16sdp_inst_769.INIT_2 = 16'h0000;
defparam ram16sdp_inst_769.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_770 (
    .DO(ram16sdp_inst_770_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_290),
    .CLK(clk)
);

defparam ram16sdp_inst_770.INIT_0 = 16'h0000;
defparam ram16sdp_inst_770.INIT_1 = 16'h0000;
defparam ram16sdp_inst_770.INIT_2 = 16'h0000;
defparam ram16sdp_inst_770.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_771 (
    .DO(ram16sdp_inst_771_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_290),
    .CLK(clk)
);

defparam ram16sdp_inst_771.INIT_0 = 16'h0000;
defparam ram16sdp_inst_771.INIT_1 = 16'h0000;
defparam ram16sdp_inst_771.INIT_2 = 16'h0000;
defparam ram16sdp_inst_771.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_772 (
    .DO(ram16sdp_inst_772_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_290),
    .CLK(clk)
);

defparam ram16sdp_inst_772.INIT_0 = 16'h0000;
defparam ram16sdp_inst_772.INIT_1 = 16'h0000;
defparam ram16sdp_inst_772.INIT_2 = 16'h0000;
defparam ram16sdp_inst_772.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_773 (
    .DO(ram16sdp_inst_773_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_290),
    .CLK(clk)
);

defparam ram16sdp_inst_773.INIT_0 = 16'h0000;
defparam ram16sdp_inst_773.INIT_1 = 16'h0000;
defparam ram16sdp_inst_773.INIT_2 = 16'h0000;
defparam ram16sdp_inst_773.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_774 (
    .DO(ram16sdp_inst_774_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_290),
    .CLK(clk)
);

defparam ram16sdp_inst_774.INIT_0 = 16'h0000;
defparam ram16sdp_inst_774.INIT_1 = 16'h0000;
defparam ram16sdp_inst_774.INIT_2 = 16'h0000;
defparam ram16sdp_inst_774.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_775 (
    .DO(ram16sdp_inst_775_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_290),
    .CLK(clk)
);

defparam ram16sdp_inst_775.INIT_0 = 16'h0000;
defparam ram16sdp_inst_775.INIT_1 = 16'h0000;
defparam ram16sdp_inst_775.INIT_2 = 16'h0000;
defparam ram16sdp_inst_775.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_776 (
    .DO(ram16sdp_inst_776_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_293),
    .CLK(clk)
);

defparam ram16sdp_inst_776.INIT_0 = 16'h0000;
defparam ram16sdp_inst_776.INIT_1 = 16'h0000;
defparam ram16sdp_inst_776.INIT_2 = 16'h0000;
defparam ram16sdp_inst_776.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_777 (
    .DO(ram16sdp_inst_777_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_293),
    .CLK(clk)
);

defparam ram16sdp_inst_777.INIT_0 = 16'h0000;
defparam ram16sdp_inst_777.INIT_1 = 16'h0000;
defparam ram16sdp_inst_777.INIT_2 = 16'h0000;
defparam ram16sdp_inst_777.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_778 (
    .DO(ram16sdp_inst_778_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_293),
    .CLK(clk)
);

defparam ram16sdp_inst_778.INIT_0 = 16'h0000;
defparam ram16sdp_inst_778.INIT_1 = 16'h0000;
defparam ram16sdp_inst_778.INIT_2 = 16'h0000;
defparam ram16sdp_inst_778.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_779 (
    .DO(ram16sdp_inst_779_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_293),
    .CLK(clk)
);

defparam ram16sdp_inst_779.INIT_0 = 16'h0000;
defparam ram16sdp_inst_779.INIT_1 = 16'h0000;
defparam ram16sdp_inst_779.INIT_2 = 16'h0000;
defparam ram16sdp_inst_779.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_780 (
    .DO(ram16sdp_inst_780_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_293),
    .CLK(clk)
);

defparam ram16sdp_inst_780.INIT_0 = 16'h0000;
defparam ram16sdp_inst_780.INIT_1 = 16'h0000;
defparam ram16sdp_inst_780.INIT_2 = 16'h0000;
defparam ram16sdp_inst_780.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_781 (
    .DO(ram16sdp_inst_781_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_293),
    .CLK(clk)
);

defparam ram16sdp_inst_781.INIT_0 = 16'h0000;
defparam ram16sdp_inst_781.INIT_1 = 16'h0000;
defparam ram16sdp_inst_781.INIT_2 = 16'h0000;
defparam ram16sdp_inst_781.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_782 (
    .DO(ram16sdp_inst_782_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_293),
    .CLK(clk)
);

defparam ram16sdp_inst_782.INIT_0 = 16'h0000;
defparam ram16sdp_inst_782.INIT_1 = 16'h0000;
defparam ram16sdp_inst_782.INIT_2 = 16'h0000;
defparam ram16sdp_inst_782.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_783 (
    .DO(ram16sdp_inst_783_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_293),
    .CLK(clk)
);

defparam ram16sdp_inst_783.INIT_0 = 16'h0000;
defparam ram16sdp_inst_783.INIT_1 = 16'h0000;
defparam ram16sdp_inst_783.INIT_2 = 16'h0000;
defparam ram16sdp_inst_783.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_784 (
    .DO(ram16sdp_inst_784_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_296),
    .CLK(clk)
);

defparam ram16sdp_inst_784.INIT_0 = 16'h0000;
defparam ram16sdp_inst_784.INIT_1 = 16'h0000;
defparam ram16sdp_inst_784.INIT_2 = 16'h0000;
defparam ram16sdp_inst_784.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_785 (
    .DO(ram16sdp_inst_785_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_296),
    .CLK(clk)
);

defparam ram16sdp_inst_785.INIT_0 = 16'h0000;
defparam ram16sdp_inst_785.INIT_1 = 16'h0000;
defparam ram16sdp_inst_785.INIT_2 = 16'h0000;
defparam ram16sdp_inst_785.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_786 (
    .DO(ram16sdp_inst_786_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_296),
    .CLK(clk)
);

defparam ram16sdp_inst_786.INIT_0 = 16'h0000;
defparam ram16sdp_inst_786.INIT_1 = 16'h0000;
defparam ram16sdp_inst_786.INIT_2 = 16'h0000;
defparam ram16sdp_inst_786.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_787 (
    .DO(ram16sdp_inst_787_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_296),
    .CLK(clk)
);

defparam ram16sdp_inst_787.INIT_0 = 16'h0000;
defparam ram16sdp_inst_787.INIT_1 = 16'h0000;
defparam ram16sdp_inst_787.INIT_2 = 16'h0000;
defparam ram16sdp_inst_787.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_788 (
    .DO(ram16sdp_inst_788_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_296),
    .CLK(clk)
);

defparam ram16sdp_inst_788.INIT_0 = 16'h0000;
defparam ram16sdp_inst_788.INIT_1 = 16'h0000;
defparam ram16sdp_inst_788.INIT_2 = 16'h0000;
defparam ram16sdp_inst_788.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_789 (
    .DO(ram16sdp_inst_789_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_296),
    .CLK(clk)
);

defparam ram16sdp_inst_789.INIT_0 = 16'h0000;
defparam ram16sdp_inst_789.INIT_1 = 16'h0000;
defparam ram16sdp_inst_789.INIT_2 = 16'h0000;
defparam ram16sdp_inst_789.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_790 (
    .DO(ram16sdp_inst_790_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_296),
    .CLK(clk)
);

defparam ram16sdp_inst_790.INIT_0 = 16'h0000;
defparam ram16sdp_inst_790.INIT_1 = 16'h0000;
defparam ram16sdp_inst_790.INIT_2 = 16'h0000;
defparam ram16sdp_inst_790.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_791 (
    .DO(ram16sdp_inst_791_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_296),
    .CLK(clk)
);

defparam ram16sdp_inst_791.INIT_0 = 16'h0000;
defparam ram16sdp_inst_791.INIT_1 = 16'h0000;
defparam ram16sdp_inst_791.INIT_2 = 16'h0000;
defparam ram16sdp_inst_791.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_792 (
    .DO(ram16sdp_inst_792_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16sdp_inst_792.INIT_0 = 16'h0000;
defparam ram16sdp_inst_792.INIT_1 = 16'h0000;
defparam ram16sdp_inst_792.INIT_2 = 16'h0000;
defparam ram16sdp_inst_792.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_793 (
    .DO(ram16sdp_inst_793_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16sdp_inst_793.INIT_0 = 16'h0000;
defparam ram16sdp_inst_793.INIT_1 = 16'h0000;
defparam ram16sdp_inst_793.INIT_2 = 16'h0000;
defparam ram16sdp_inst_793.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_794 (
    .DO(ram16sdp_inst_794_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16sdp_inst_794.INIT_0 = 16'h0000;
defparam ram16sdp_inst_794.INIT_1 = 16'h0000;
defparam ram16sdp_inst_794.INIT_2 = 16'h0000;
defparam ram16sdp_inst_794.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_795 (
    .DO(ram16sdp_inst_795_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16sdp_inst_795.INIT_0 = 16'h0000;
defparam ram16sdp_inst_795.INIT_1 = 16'h0000;
defparam ram16sdp_inst_795.INIT_2 = 16'h0000;
defparam ram16sdp_inst_795.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_796 (
    .DO(ram16sdp_inst_796_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16sdp_inst_796.INIT_0 = 16'h0000;
defparam ram16sdp_inst_796.INIT_1 = 16'h0000;
defparam ram16sdp_inst_796.INIT_2 = 16'h0000;
defparam ram16sdp_inst_796.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_797 (
    .DO(ram16sdp_inst_797_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16sdp_inst_797.INIT_0 = 16'h0000;
defparam ram16sdp_inst_797.INIT_1 = 16'h0000;
defparam ram16sdp_inst_797.INIT_2 = 16'h0000;
defparam ram16sdp_inst_797.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_798 (
    .DO(ram16sdp_inst_798_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16sdp_inst_798.INIT_0 = 16'h0000;
defparam ram16sdp_inst_798.INIT_1 = 16'h0000;
defparam ram16sdp_inst_798.INIT_2 = 16'h0000;
defparam ram16sdp_inst_798.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_799 (
    .DO(ram16sdp_inst_799_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16sdp_inst_799.INIT_0 = 16'h0000;
defparam ram16sdp_inst_799.INIT_1 = 16'h0000;
defparam ram16sdp_inst_799.INIT_2 = 16'h0000;
defparam ram16sdp_inst_799.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_800 (
    .DO(ram16sdp_inst_800_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_302),
    .CLK(clk)
);

defparam ram16sdp_inst_800.INIT_0 = 16'h0000;
defparam ram16sdp_inst_800.INIT_1 = 16'h0000;
defparam ram16sdp_inst_800.INIT_2 = 16'h0000;
defparam ram16sdp_inst_800.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_801 (
    .DO(ram16sdp_inst_801_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_302),
    .CLK(clk)
);

defparam ram16sdp_inst_801.INIT_0 = 16'h0000;
defparam ram16sdp_inst_801.INIT_1 = 16'h0000;
defparam ram16sdp_inst_801.INIT_2 = 16'h0000;
defparam ram16sdp_inst_801.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_802 (
    .DO(ram16sdp_inst_802_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_302),
    .CLK(clk)
);

defparam ram16sdp_inst_802.INIT_0 = 16'h0000;
defparam ram16sdp_inst_802.INIT_1 = 16'h0000;
defparam ram16sdp_inst_802.INIT_2 = 16'h0000;
defparam ram16sdp_inst_802.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_803 (
    .DO(ram16sdp_inst_803_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_302),
    .CLK(clk)
);

defparam ram16sdp_inst_803.INIT_0 = 16'h0000;
defparam ram16sdp_inst_803.INIT_1 = 16'h0000;
defparam ram16sdp_inst_803.INIT_2 = 16'h0000;
defparam ram16sdp_inst_803.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_804 (
    .DO(ram16sdp_inst_804_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_302),
    .CLK(clk)
);

defparam ram16sdp_inst_804.INIT_0 = 16'h0000;
defparam ram16sdp_inst_804.INIT_1 = 16'h0000;
defparam ram16sdp_inst_804.INIT_2 = 16'h0000;
defparam ram16sdp_inst_804.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_805 (
    .DO(ram16sdp_inst_805_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_302),
    .CLK(clk)
);

defparam ram16sdp_inst_805.INIT_0 = 16'h0000;
defparam ram16sdp_inst_805.INIT_1 = 16'h0000;
defparam ram16sdp_inst_805.INIT_2 = 16'h0000;
defparam ram16sdp_inst_805.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_806 (
    .DO(ram16sdp_inst_806_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_302),
    .CLK(clk)
);

defparam ram16sdp_inst_806.INIT_0 = 16'h0000;
defparam ram16sdp_inst_806.INIT_1 = 16'h0000;
defparam ram16sdp_inst_806.INIT_2 = 16'h0000;
defparam ram16sdp_inst_806.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_807 (
    .DO(ram16sdp_inst_807_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_302),
    .CLK(clk)
);

defparam ram16sdp_inst_807.INIT_0 = 16'h0000;
defparam ram16sdp_inst_807.INIT_1 = 16'h0000;
defparam ram16sdp_inst_807.INIT_2 = 16'h0000;
defparam ram16sdp_inst_807.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_808 (
    .DO(ram16sdp_inst_808_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_305),
    .CLK(clk)
);

defparam ram16sdp_inst_808.INIT_0 = 16'h0000;
defparam ram16sdp_inst_808.INIT_1 = 16'h0000;
defparam ram16sdp_inst_808.INIT_2 = 16'h0000;
defparam ram16sdp_inst_808.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_809 (
    .DO(ram16sdp_inst_809_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_305),
    .CLK(clk)
);

defparam ram16sdp_inst_809.INIT_0 = 16'h0000;
defparam ram16sdp_inst_809.INIT_1 = 16'h0000;
defparam ram16sdp_inst_809.INIT_2 = 16'h0000;
defparam ram16sdp_inst_809.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_810 (
    .DO(ram16sdp_inst_810_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_305),
    .CLK(clk)
);

defparam ram16sdp_inst_810.INIT_0 = 16'h0000;
defparam ram16sdp_inst_810.INIT_1 = 16'h0000;
defparam ram16sdp_inst_810.INIT_2 = 16'h0000;
defparam ram16sdp_inst_810.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_811 (
    .DO(ram16sdp_inst_811_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_305),
    .CLK(clk)
);

defparam ram16sdp_inst_811.INIT_0 = 16'h0000;
defparam ram16sdp_inst_811.INIT_1 = 16'h0000;
defparam ram16sdp_inst_811.INIT_2 = 16'h0000;
defparam ram16sdp_inst_811.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_812 (
    .DO(ram16sdp_inst_812_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_305),
    .CLK(clk)
);

defparam ram16sdp_inst_812.INIT_0 = 16'h0000;
defparam ram16sdp_inst_812.INIT_1 = 16'h0000;
defparam ram16sdp_inst_812.INIT_2 = 16'h0000;
defparam ram16sdp_inst_812.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_813 (
    .DO(ram16sdp_inst_813_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_305),
    .CLK(clk)
);

defparam ram16sdp_inst_813.INIT_0 = 16'h0000;
defparam ram16sdp_inst_813.INIT_1 = 16'h0000;
defparam ram16sdp_inst_813.INIT_2 = 16'h0000;
defparam ram16sdp_inst_813.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_814 (
    .DO(ram16sdp_inst_814_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_305),
    .CLK(clk)
);

defparam ram16sdp_inst_814.INIT_0 = 16'h0000;
defparam ram16sdp_inst_814.INIT_1 = 16'h0000;
defparam ram16sdp_inst_814.INIT_2 = 16'h0000;
defparam ram16sdp_inst_814.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_815 (
    .DO(ram16sdp_inst_815_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_305),
    .CLK(clk)
);

defparam ram16sdp_inst_815.INIT_0 = 16'h0000;
defparam ram16sdp_inst_815.INIT_1 = 16'h0000;
defparam ram16sdp_inst_815.INIT_2 = 16'h0000;
defparam ram16sdp_inst_815.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_816 (
    .DO(ram16sdp_inst_816_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_308),
    .CLK(clk)
);

defparam ram16sdp_inst_816.INIT_0 = 16'h0000;
defparam ram16sdp_inst_816.INIT_1 = 16'h0000;
defparam ram16sdp_inst_816.INIT_2 = 16'h0000;
defparam ram16sdp_inst_816.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_817 (
    .DO(ram16sdp_inst_817_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_308),
    .CLK(clk)
);

defparam ram16sdp_inst_817.INIT_0 = 16'h0000;
defparam ram16sdp_inst_817.INIT_1 = 16'h0000;
defparam ram16sdp_inst_817.INIT_2 = 16'h0000;
defparam ram16sdp_inst_817.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_818 (
    .DO(ram16sdp_inst_818_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_308),
    .CLK(clk)
);

defparam ram16sdp_inst_818.INIT_0 = 16'h0000;
defparam ram16sdp_inst_818.INIT_1 = 16'h0000;
defparam ram16sdp_inst_818.INIT_2 = 16'h0000;
defparam ram16sdp_inst_818.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_819 (
    .DO(ram16sdp_inst_819_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_308),
    .CLK(clk)
);

defparam ram16sdp_inst_819.INIT_0 = 16'h0000;
defparam ram16sdp_inst_819.INIT_1 = 16'h0000;
defparam ram16sdp_inst_819.INIT_2 = 16'h0000;
defparam ram16sdp_inst_819.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_820 (
    .DO(ram16sdp_inst_820_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_308),
    .CLK(clk)
);

defparam ram16sdp_inst_820.INIT_0 = 16'h0000;
defparam ram16sdp_inst_820.INIT_1 = 16'h0000;
defparam ram16sdp_inst_820.INIT_2 = 16'h0000;
defparam ram16sdp_inst_820.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_821 (
    .DO(ram16sdp_inst_821_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_308),
    .CLK(clk)
);

defparam ram16sdp_inst_821.INIT_0 = 16'h0000;
defparam ram16sdp_inst_821.INIT_1 = 16'h0000;
defparam ram16sdp_inst_821.INIT_2 = 16'h0000;
defparam ram16sdp_inst_821.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_822 (
    .DO(ram16sdp_inst_822_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_308),
    .CLK(clk)
);

defparam ram16sdp_inst_822.INIT_0 = 16'h0000;
defparam ram16sdp_inst_822.INIT_1 = 16'h0000;
defparam ram16sdp_inst_822.INIT_2 = 16'h0000;
defparam ram16sdp_inst_822.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_823 (
    .DO(ram16sdp_inst_823_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_308),
    .CLK(clk)
);

defparam ram16sdp_inst_823.INIT_0 = 16'h0000;
defparam ram16sdp_inst_823.INIT_1 = 16'h0000;
defparam ram16sdp_inst_823.INIT_2 = 16'h0000;
defparam ram16sdp_inst_823.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_824 (
    .DO(ram16sdp_inst_824_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16sdp_inst_824.INIT_0 = 16'h0000;
defparam ram16sdp_inst_824.INIT_1 = 16'h0000;
defparam ram16sdp_inst_824.INIT_2 = 16'h0000;
defparam ram16sdp_inst_824.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_825 (
    .DO(ram16sdp_inst_825_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16sdp_inst_825.INIT_0 = 16'h0000;
defparam ram16sdp_inst_825.INIT_1 = 16'h0000;
defparam ram16sdp_inst_825.INIT_2 = 16'h0000;
defparam ram16sdp_inst_825.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_826 (
    .DO(ram16sdp_inst_826_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16sdp_inst_826.INIT_0 = 16'h0000;
defparam ram16sdp_inst_826.INIT_1 = 16'h0000;
defparam ram16sdp_inst_826.INIT_2 = 16'h0000;
defparam ram16sdp_inst_826.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_827 (
    .DO(ram16sdp_inst_827_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16sdp_inst_827.INIT_0 = 16'h0000;
defparam ram16sdp_inst_827.INIT_1 = 16'h0000;
defparam ram16sdp_inst_827.INIT_2 = 16'h0000;
defparam ram16sdp_inst_827.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_828 (
    .DO(ram16sdp_inst_828_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16sdp_inst_828.INIT_0 = 16'h0000;
defparam ram16sdp_inst_828.INIT_1 = 16'h0000;
defparam ram16sdp_inst_828.INIT_2 = 16'h0000;
defparam ram16sdp_inst_828.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_829 (
    .DO(ram16sdp_inst_829_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16sdp_inst_829.INIT_0 = 16'h0000;
defparam ram16sdp_inst_829.INIT_1 = 16'h0000;
defparam ram16sdp_inst_829.INIT_2 = 16'h0000;
defparam ram16sdp_inst_829.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_830 (
    .DO(ram16sdp_inst_830_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16sdp_inst_830.INIT_0 = 16'h0000;
defparam ram16sdp_inst_830.INIT_1 = 16'h0000;
defparam ram16sdp_inst_830.INIT_2 = 16'h0000;
defparam ram16sdp_inst_830.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_831 (
    .DO(ram16sdp_inst_831_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16sdp_inst_831.INIT_0 = 16'h0000;
defparam ram16sdp_inst_831.INIT_1 = 16'h0000;
defparam ram16sdp_inst_831.INIT_2 = 16'h0000;
defparam ram16sdp_inst_831.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_832 (
    .DO(ram16sdp_inst_832_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_314),
    .CLK(clk)
);

defparam ram16sdp_inst_832.INIT_0 = 16'h0000;
defparam ram16sdp_inst_832.INIT_1 = 16'h0000;
defparam ram16sdp_inst_832.INIT_2 = 16'h0000;
defparam ram16sdp_inst_832.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_833 (
    .DO(ram16sdp_inst_833_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_314),
    .CLK(clk)
);

defparam ram16sdp_inst_833.INIT_0 = 16'h0000;
defparam ram16sdp_inst_833.INIT_1 = 16'h0000;
defparam ram16sdp_inst_833.INIT_2 = 16'h0000;
defparam ram16sdp_inst_833.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_834 (
    .DO(ram16sdp_inst_834_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_314),
    .CLK(clk)
);

defparam ram16sdp_inst_834.INIT_0 = 16'h0000;
defparam ram16sdp_inst_834.INIT_1 = 16'h0000;
defparam ram16sdp_inst_834.INIT_2 = 16'h0000;
defparam ram16sdp_inst_834.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_835 (
    .DO(ram16sdp_inst_835_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_314),
    .CLK(clk)
);

defparam ram16sdp_inst_835.INIT_0 = 16'h0000;
defparam ram16sdp_inst_835.INIT_1 = 16'h0000;
defparam ram16sdp_inst_835.INIT_2 = 16'h0000;
defparam ram16sdp_inst_835.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_836 (
    .DO(ram16sdp_inst_836_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_314),
    .CLK(clk)
);

defparam ram16sdp_inst_836.INIT_0 = 16'h0000;
defparam ram16sdp_inst_836.INIT_1 = 16'h0000;
defparam ram16sdp_inst_836.INIT_2 = 16'h0000;
defparam ram16sdp_inst_836.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_837 (
    .DO(ram16sdp_inst_837_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_314),
    .CLK(clk)
);

defparam ram16sdp_inst_837.INIT_0 = 16'h0000;
defparam ram16sdp_inst_837.INIT_1 = 16'h0000;
defparam ram16sdp_inst_837.INIT_2 = 16'h0000;
defparam ram16sdp_inst_837.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_838 (
    .DO(ram16sdp_inst_838_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_314),
    .CLK(clk)
);

defparam ram16sdp_inst_838.INIT_0 = 16'h0000;
defparam ram16sdp_inst_838.INIT_1 = 16'h0000;
defparam ram16sdp_inst_838.INIT_2 = 16'h0000;
defparam ram16sdp_inst_838.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_839 (
    .DO(ram16sdp_inst_839_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_314),
    .CLK(clk)
);

defparam ram16sdp_inst_839.INIT_0 = 16'h0000;
defparam ram16sdp_inst_839.INIT_1 = 16'h0000;
defparam ram16sdp_inst_839.INIT_2 = 16'h0000;
defparam ram16sdp_inst_839.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_840 (
    .DO(ram16sdp_inst_840_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_317),
    .CLK(clk)
);

defparam ram16sdp_inst_840.INIT_0 = 16'h0000;
defparam ram16sdp_inst_840.INIT_1 = 16'h0000;
defparam ram16sdp_inst_840.INIT_2 = 16'h0000;
defparam ram16sdp_inst_840.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_841 (
    .DO(ram16sdp_inst_841_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_317),
    .CLK(clk)
);

defparam ram16sdp_inst_841.INIT_0 = 16'h0000;
defparam ram16sdp_inst_841.INIT_1 = 16'h0000;
defparam ram16sdp_inst_841.INIT_2 = 16'h0000;
defparam ram16sdp_inst_841.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_842 (
    .DO(ram16sdp_inst_842_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_317),
    .CLK(clk)
);

defparam ram16sdp_inst_842.INIT_0 = 16'h0000;
defparam ram16sdp_inst_842.INIT_1 = 16'h0000;
defparam ram16sdp_inst_842.INIT_2 = 16'h0000;
defparam ram16sdp_inst_842.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_843 (
    .DO(ram16sdp_inst_843_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_317),
    .CLK(clk)
);

defparam ram16sdp_inst_843.INIT_0 = 16'h0000;
defparam ram16sdp_inst_843.INIT_1 = 16'h0000;
defparam ram16sdp_inst_843.INIT_2 = 16'h0000;
defparam ram16sdp_inst_843.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_844 (
    .DO(ram16sdp_inst_844_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_317),
    .CLK(clk)
);

defparam ram16sdp_inst_844.INIT_0 = 16'h0000;
defparam ram16sdp_inst_844.INIT_1 = 16'h0000;
defparam ram16sdp_inst_844.INIT_2 = 16'h0000;
defparam ram16sdp_inst_844.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_845 (
    .DO(ram16sdp_inst_845_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_317),
    .CLK(clk)
);

defparam ram16sdp_inst_845.INIT_0 = 16'h0000;
defparam ram16sdp_inst_845.INIT_1 = 16'h0000;
defparam ram16sdp_inst_845.INIT_2 = 16'h0000;
defparam ram16sdp_inst_845.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_846 (
    .DO(ram16sdp_inst_846_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_317),
    .CLK(clk)
);

defparam ram16sdp_inst_846.INIT_0 = 16'h0000;
defparam ram16sdp_inst_846.INIT_1 = 16'h0000;
defparam ram16sdp_inst_846.INIT_2 = 16'h0000;
defparam ram16sdp_inst_846.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_847 (
    .DO(ram16sdp_inst_847_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_317),
    .CLK(clk)
);

defparam ram16sdp_inst_847.INIT_0 = 16'h0000;
defparam ram16sdp_inst_847.INIT_1 = 16'h0000;
defparam ram16sdp_inst_847.INIT_2 = 16'h0000;
defparam ram16sdp_inst_847.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_848 (
    .DO(ram16sdp_inst_848_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_320),
    .CLK(clk)
);

defparam ram16sdp_inst_848.INIT_0 = 16'h0000;
defparam ram16sdp_inst_848.INIT_1 = 16'h0000;
defparam ram16sdp_inst_848.INIT_2 = 16'h0000;
defparam ram16sdp_inst_848.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_849 (
    .DO(ram16sdp_inst_849_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_320),
    .CLK(clk)
);

defparam ram16sdp_inst_849.INIT_0 = 16'h0000;
defparam ram16sdp_inst_849.INIT_1 = 16'h0000;
defparam ram16sdp_inst_849.INIT_2 = 16'h0000;
defparam ram16sdp_inst_849.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_850 (
    .DO(ram16sdp_inst_850_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_320),
    .CLK(clk)
);

defparam ram16sdp_inst_850.INIT_0 = 16'h0000;
defparam ram16sdp_inst_850.INIT_1 = 16'h0000;
defparam ram16sdp_inst_850.INIT_2 = 16'h0000;
defparam ram16sdp_inst_850.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_851 (
    .DO(ram16sdp_inst_851_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_320),
    .CLK(clk)
);

defparam ram16sdp_inst_851.INIT_0 = 16'h0000;
defparam ram16sdp_inst_851.INIT_1 = 16'h0000;
defparam ram16sdp_inst_851.INIT_2 = 16'h0000;
defparam ram16sdp_inst_851.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_852 (
    .DO(ram16sdp_inst_852_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_320),
    .CLK(clk)
);

defparam ram16sdp_inst_852.INIT_0 = 16'h0000;
defparam ram16sdp_inst_852.INIT_1 = 16'h0000;
defparam ram16sdp_inst_852.INIT_2 = 16'h0000;
defparam ram16sdp_inst_852.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_853 (
    .DO(ram16sdp_inst_853_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_320),
    .CLK(clk)
);

defparam ram16sdp_inst_853.INIT_0 = 16'h0000;
defparam ram16sdp_inst_853.INIT_1 = 16'h0000;
defparam ram16sdp_inst_853.INIT_2 = 16'h0000;
defparam ram16sdp_inst_853.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_854 (
    .DO(ram16sdp_inst_854_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_320),
    .CLK(clk)
);

defparam ram16sdp_inst_854.INIT_0 = 16'h0000;
defparam ram16sdp_inst_854.INIT_1 = 16'h0000;
defparam ram16sdp_inst_854.INIT_2 = 16'h0000;
defparam ram16sdp_inst_854.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_855 (
    .DO(ram16sdp_inst_855_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_320),
    .CLK(clk)
);

defparam ram16sdp_inst_855.INIT_0 = 16'h0000;
defparam ram16sdp_inst_855.INIT_1 = 16'h0000;
defparam ram16sdp_inst_855.INIT_2 = 16'h0000;
defparam ram16sdp_inst_855.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_856 (
    .DO(ram16sdp_inst_856_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16sdp_inst_856.INIT_0 = 16'h0000;
defparam ram16sdp_inst_856.INIT_1 = 16'h0000;
defparam ram16sdp_inst_856.INIT_2 = 16'h0000;
defparam ram16sdp_inst_856.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_857 (
    .DO(ram16sdp_inst_857_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16sdp_inst_857.INIT_0 = 16'h0000;
defparam ram16sdp_inst_857.INIT_1 = 16'h0000;
defparam ram16sdp_inst_857.INIT_2 = 16'h0000;
defparam ram16sdp_inst_857.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_858 (
    .DO(ram16sdp_inst_858_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16sdp_inst_858.INIT_0 = 16'h0000;
defparam ram16sdp_inst_858.INIT_1 = 16'h0000;
defparam ram16sdp_inst_858.INIT_2 = 16'h0000;
defparam ram16sdp_inst_858.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_859 (
    .DO(ram16sdp_inst_859_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16sdp_inst_859.INIT_0 = 16'h0000;
defparam ram16sdp_inst_859.INIT_1 = 16'h0000;
defparam ram16sdp_inst_859.INIT_2 = 16'h0000;
defparam ram16sdp_inst_859.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_860 (
    .DO(ram16sdp_inst_860_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16sdp_inst_860.INIT_0 = 16'h0000;
defparam ram16sdp_inst_860.INIT_1 = 16'h0000;
defparam ram16sdp_inst_860.INIT_2 = 16'h0000;
defparam ram16sdp_inst_860.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_861 (
    .DO(ram16sdp_inst_861_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16sdp_inst_861.INIT_0 = 16'h0000;
defparam ram16sdp_inst_861.INIT_1 = 16'h0000;
defparam ram16sdp_inst_861.INIT_2 = 16'h0000;
defparam ram16sdp_inst_861.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_862 (
    .DO(ram16sdp_inst_862_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16sdp_inst_862.INIT_0 = 16'h0000;
defparam ram16sdp_inst_862.INIT_1 = 16'h0000;
defparam ram16sdp_inst_862.INIT_2 = 16'h0000;
defparam ram16sdp_inst_862.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_863 (
    .DO(ram16sdp_inst_863_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16sdp_inst_863.INIT_0 = 16'h0000;
defparam ram16sdp_inst_863.INIT_1 = 16'h0000;
defparam ram16sdp_inst_863.INIT_2 = 16'h0000;
defparam ram16sdp_inst_863.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_864 (
    .DO(ram16sdp_inst_864_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_326),
    .CLK(clk)
);

defparam ram16sdp_inst_864.INIT_0 = 16'h0000;
defparam ram16sdp_inst_864.INIT_1 = 16'h0000;
defparam ram16sdp_inst_864.INIT_2 = 16'h0000;
defparam ram16sdp_inst_864.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_865 (
    .DO(ram16sdp_inst_865_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_326),
    .CLK(clk)
);

defparam ram16sdp_inst_865.INIT_0 = 16'h0000;
defparam ram16sdp_inst_865.INIT_1 = 16'h0000;
defparam ram16sdp_inst_865.INIT_2 = 16'h0000;
defparam ram16sdp_inst_865.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_866 (
    .DO(ram16sdp_inst_866_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_326),
    .CLK(clk)
);

defparam ram16sdp_inst_866.INIT_0 = 16'h0000;
defparam ram16sdp_inst_866.INIT_1 = 16'h0000;
defparam ram16sdp_inst_866.INIT_2 = 16'h0000;
defparam ram16sdp_inst_866.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_867 (
    .DO(ram16sdp_inst_867_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_326),
    .CLK(clk)
);

defparam ram16sdp_inst_867.INIT_0 = 16'h0000;
defparam ram16sdp_inst_867.INIT_1 = 16'h0000;
defparam ram16sdp_inst_867.INIT_2 = 16'h0000;
defparam ram16sdp_inst_867.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_868 (
    .DO(ram16sdp_inst_868_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_326),
    .CLK(clk)
);

defparam ram16sdp_inst_868.INIT_0 = 16'h0000;
defparam ram16sdp_inst_868.INIT_1 = 16'h0000;
defparam ram16sdp_inst_868.INIT_2 = 16'h0000;
defparam ram16sdp_inst_868.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_869 (
    .DO(ram16sdp_inst_869_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_326),
    .CLK(clk)
);

defparam ram16sdp_inst_869.INIT_0 = 16'h0000;
defparam ram16sdp_inst_869.INIT_1 = 16'h0000;
defparam ram16sdp_inst_869.INIT_2 = 16'h0000;
defparam ram16sdp_inst_869.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_870 (
    .DO(ram16sdp_inst_870_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_326),
    .CLK(clk)
);

defparam ram16sdp_inst_870.INIT_0 = 16'h0000;
defparam ram16sdp_inst_870.INIT_1 = 16'h0000;
defparam ram16sdp_inst_870.INIT_2 = 16'h0000;
defparam ram16sdp_inst_870.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_871 (
    .DO(ram16sdp_inst_871_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_326),
    .CLK(clk)
);

defparam ram16sdp_inst_871.INIT_0 = 16'h0000;
defparam ram16sdp_inst_871.INIT_1 = 16'h0000;
defparam ram16sdp_inst_871.INIT_2 = 16'h0000;
defparam ram16sdp_inst_871.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_872 (
    .DO(ram16sdp_inst_872_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_329),
    .CLK(clk)
);

defparam ram16sdp_inst_872.INIT_0 = 16'h0000;
defparam ram16sdp_inst_872.INIT_1 = 16'h0000;
defparam ram16sdp_inst_872.INIT_2 = 16'h0000;
defparam ram16sdp_inst_872.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_873 (
    .DO(ram16sdp_inst_873_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_329),
    .CLK(clk)
);

defparam ram16sdp_inst_873.INIT_0 = 16'h0000;
defparam ram16sdp_inst_873.INIT_1 = 16'h0000;
defparam ram16sdp_inst_873.INIT_2 = 16'h0000;
defparam ram16sdp_inst_873.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_874 (
    .DO(ram16sdp_inst_874_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_329),
    .CLK(clk)
);

defparam ram16sdp_inst_874.INIT_0 = 16'h0000;
defparam ram16sdp_inst_874.INIT_1 = 16'h0000;
defparam ram16sdp_inst_874.INIT_2 = 16'h0000;
defparam ram16sdp_inst_874.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_875 (
    .DO(ram16sdp_inst_875_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_329),
    .CLK(clk)
);

defparam ram16sdp_inst_875.INIT_0 = 16'h0000;
defparam ram16sdp_inst_875.INIT_1 = 16'h0000;
defparam ram16sdp_inst_875.INIT_2 = 16'h0000;
defparam ram16sdp_inst_875.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_876 (
    .DO(ram16sdp_inst_876_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_329),
    .CLK(clk)
);

defparam ram16sdp_inst_876.INIT_0 = 16'h0000;
defparam ram16sdp_inst_876.INIT_1 = 16'h0000;
defparam ram16sdp_inst_876.INIT_2 = 16'h0000;
defparam ram16sdp_inst_876.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_877 (
    .DO(ram16sdp_inst_877_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_329),
    .CLK(clk)
);

defparam ram16sdp_inst_877.INIT_0 = 16'h0000;
defparam ram16sdp_inst_877.INIT_1 = 16'h0000;
defparam ram16sdp_inst_877.INIT_2 = 16'h0000;
defparam ram16sdp_inst_877.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_878 (
    .DO(ram16sdp_inst_878_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_329),
    .CLK(clk)
);

defparam ram16sdp_inst_878.INIT_0 = 16'h0000;
defparam ram16sdp_inst_878.INIT_1 = 16'h0000;
defparam ram16sdp_inst_878.INIT_2 = 16'h0000;
defparam ram16sdp_inst_878.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_879 (
    .DO(ram16sdp_inst_879_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_329),
    .CLK(clk)
);

defparam ram16sdp_inst_879.INIT_0 = 16'h0000;
defparam ram16sdp_inst_879.INIT_1 = 16'h0000;
defparam ram16sdp_inst_879.INIT_2 = 16'h0000;
defparam ram16sdp_inst_879.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_880 (
    .DO(ram16sdp_inst_880_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_332),
    .CLK(clk)
);

defparam ram16sdp_inst_880.INIT_0 = 16'h0000;
defparam ram16sdp_inst_880.INIT_1 = 16'h0000;
defparam ram16sdp_inst_880.INIT_2 = 16'h0000;
defparam ram16sdp_inst_880.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_881 (
    .DO(ram16sdp_inst_881_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_332),
    .CLK(clk)
);

defparam ram16sdp_inst_881.INIT_0 = 16'h0000;
defparam ram16sdp_inst_881.INIT_1 = 16'h0000;
defparam ram16sdp_inst_881.INIT_2 = 16'h0000;
defparam ram16sdp_inst_881.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_882 (
    .DO(ram16sdp_inst_882_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_332),
    .CLK(clk)
);

defparam ram16sdp_inst_882.INIT_0 = 16'h0000;
defparam ram16sdp_inst_882.INIT_1 = 16'h0000;
defparam ram16sdp_inst_882.INIT_2 = 16'h0000;
defparam ram16sdp_inst_882.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_883 (
    .DO(ram16sdp_inst_883_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_332),
    .CLK(clk)
);

defparam ram16sdp_inst_883.INIT_0 = 16'h0000;
defparam ram16sdp_inst_883.INIT_1 = 16'h0000;
defparam ram16sdp_inst_883.INIT_2 = 16'h0000;
defparam ram16sdp_inst_883.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_884 (
    .DO(ram16sdp_inst_884_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_332),
    .CLK(clk)
);

defparam ram16sdp_inst_884.INIT_0 = 16'h0000;
defparam ram16sdp_inst_884.INIT_1 = 16'h0000;
defparam ram16sdp_inst_884.INIT_2 = 16'h0000;
defparam ram16sdp_inst_884.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_885 (
    .DO(ram16sdp_inst_885_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_332),
    .CLK(clk)
);

defparam ram16sdp_inst_885.INIT_0 = 16'h0000;
defparam ram16sdp_inst_885.INIT_1 = 16'h0000;
defparam ram16sdp_inst_885.INIT_2 = 16'h0000;
defparam ram16sdp_inst_885.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_886 (
    .DO(ram16sdp_inst_886_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_332),
    .CLK(clk)
);

defparam ram16sdp_inst_886.INIT_0 = 16'h0000;
defparam ram16sdp_inst_886.INIT_1 = 16'h0000;
defparam ram16sdp_inst_886.INIT_2 = 16'h0000;
defparam ram16sdp_inst_886.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_887 (
    .DO(ram16sdp_inst_887_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_332),
    .CLK(clk)
);

defparam ram16sdp_inst_887.INIT_0 = 16'h0000;
defparam ram16sdp_inst_887.INIT_1 = 16'h0000;
defparam ram16sdp_inst_887.INIT_2 = 16'h0000;
defparam ram16sdp_inst_887.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_888 (
    .DO(ram16sdp_inst_888_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16sdp_inst_888.INIT_0 = 16'h0000;
defparam ram16sdp_inst_888.INIT_1 = 16'h0000;
defparam ram16sdp_inst_888.INIT_2 = 16'h0000;
defparam ram16sdp_inst_888.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_889 (
    .DO(ram16sdp_inst_889_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16sdp_inst_889.INIT_0 = 16'h0000;
defparam ram16sdp_inst_889.INIT_1 = 16'h0000;
defparam ram16sdp_inst_889.INIT_2 = 16'h0000;
defparam ram16sdp_inst_889.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_890 (
    .DO(ram16sdp_inst_890_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16sdp_inst_890.INIT_0 = 16'h0000;
defparam ram16sdp_inst_890.INIT_1 = 16'h0000;
defparam ram16sdp_inst_890.INIT_2 = 16'h0000;
defparam ram16sdp_inst_890.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_891 (
    .DO(ram16sdp_inst_891_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16sdp_inst_891.INIT_0 = 16'h0000;
defparam ram16sdp_inst_891.INIT_1 = 16'h0000;
defparam ram16sdp_inst_891.INIT_2 = 16'h0000;
defparam ram16sdp_inst_891.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_892 (
    .DO(ram16sdp_inst_892_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16sdp_inst_892.INIT_0 = 16'h0000;
defparam ram16sdp_inst_892.INIT_1 = 16'h0000;
defparam ram16sdp_inst_892.INIT_2 = 16'h0000;
defparam ram16sdp_inst_892.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_893 (
    .DO(ram16sdp_inst_893_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16sdp_inst_893.INIT_0 = 16'h0000;
defparam ram16sdp_inst_893.INIT_1 = 16'h0000;
defparam ram16sdp_inst_893.INIT_2 = 16'h0000;
defparam ram16sdp_inst_893.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_894 (
    .DO(ram16sdp_inst_894_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16sdp_inst_894.INIT_0 = 16'h0000;
defparam ram16sdp_inst_894.INIT_1 = 16'h0000;
defparam ram16sdp_inst_894.INIT_2 = 16'h0000;
defparam ram16sdp_inst_894.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_895 (
    .DO(ram16sdp_inst_895_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16sdp_inst_895.INIT_0 = 16'h0000;
defparam ram16sdp_inst_895.INIT_1 = 16'h0000;
defparam ram16sdp_inst_895.INIT_2 = 16'h0000;
defparam ram16sdp_inst_895.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_896 (
    .DO(ram16sdp_inst_896_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_338),
    .CLK(clk)
);

defparam ram16sdp_inst_896.INIT_0 = 16'h0000;
defparam ram16sdp_inst_896.INIT_1 = 16'h0000;
defparam ram16sdp_inst_896.INIT_2 = 16'h0000;
defparam ram16sdp_inst_896.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_897 (
    .DO(ram16sdp_inst_897_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_338),
    .CLK(clk)
);

defparam ram16sdp_inst_897.INIT_0 = 16'h0000;
defparam ram16sdp_inst_897.INIT_1 = 16'h0000;
defparam ram16sdp_inst_897.INIT_2 = 16'h0000;
defparam ram16sdp_inst_897.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_898 (
    .DO(ram16sdp_inst_898_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_338),
    .CLK(clk)
);

defparam ram16sdp_inst_898.INIT_0 = 16'h0000;
defparam ram16sdp_inst_898.INIT_1 = 16'h0000;
defparam ram16sdp_inst_898.INIT_2 = 16'h0000;
defparam ram16sdp_inst_898.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_899 (
    .DO(ram16sdp_inst_899_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_338),
    .CLK(clk)
);

defparam ram16sdp_inst_899.INIT_0 = 16'h0000;
defparam ram16sdp_inst_899.INIT_1 = 16'h0000;
defparam ram16sdp_inst_899.INIT_2 = 16'h0000;
defparam ram16sdp_inst_899.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_900 (
    .DO(ram16sdp_inst_900_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_338),
    .CLK(clk)
);

defparam ram16sdp_inst_900.INIT_0 = 16'h0000;
defparam ram16sdp_inst_900.INIT_1 = 16'h0000;
defparam ram16sdp_inst_900.INIT_2 = 16'h0000;
defparam ram16sdp_inst_900.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_901 (
    .DO(ram16sdp_inst_901_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_338),
    .CLK(clk)
);

defparam ram16sdp_inst_901.INIT_0 = 16'h0000;
defparam ram16sdp_inst_901.INIT_1 = 16'h0000;
defparam ram16sdp_inst_901.INIT_2 = 16'h0000;
defparam ram16sdp_inst_901.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_902 (
    .DO(ram16sdp_inst_902_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_338),
    .CLK(clk)
);

defparam ram16sdp_inst_902.INIT_0 = 16'h0000;
defparam ram16sdp_inst_902.INIT_1 = 16'h0000;
defparam ram16sdp_inst_902.INIT_2 = 16'h0000;
defparam ram16sdp_inst_902.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_903 (
    .DO(ram16sdp_inst_903_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_338),
    .CLK(clk)
);

defparam ram16sdp_inst_903.INIT_0 = 16'h0000;
defparam ram16sdp_inst_903.INIT_1 = 16'h0000;
defparam ram16sdp_inst_903.INIT_2 = 16'h0000;
defparam ram16sdp_inst_903.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_904 (
    .DO(ram16sdp_inst_904_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_341),
    .CLK(clk)
);

defparam ram16sdp_inst_904.INIT_0 = 16'h0000;
defparam ram16sdp_inst_904.INIT_1 = 16'h0000;
defparam ram16sdp_inst_904.INIT_2 = 16'h0000;
defparam ram16sdp_inst_904.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_905 (
    .DO(ram16sdp_inst_905_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_341),
    .CLK(clk)
);

defparam ram16sdp_inst_905.INIT_0 = 16'h0000;
defparam ram16sdp_inst_905.INIT_1 = 16'h0000;
defparam ram16sdp_inst_905.INIT_2 = 16'h0000;
defparam ram16sdp_inst_905.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_906 (
    .DO(ram16sdp_inst_906_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_341),
    .CLK(clk)
);

defparam ram16sdp_inst_906.INIT_0 = 16'h0000;
defparam ram16sdp_inst_906.INIT_1 = 16'h0000;
defparam ram16sdp_inst_906.INIT_2 = 16'h0000;
defparam ram16sdp_inst_906.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_907 (
    .DO(ram16sdp_inst_907_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_341),
    .CLK(clk)
);

defparam ram16sdp_inst_907.INIT_0 = 16'h0000;
defparam ram16sdp_inst_907.INIT_1 = 16'h0000;
defparam ram16sdp_inst_907.INIT_2 = 16'h0000;
defparam ram16sdp_inst_907.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_908 (
    .DO(ram16sdp_inst_908_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_341),
    .CLK(clk)
);

defparam ram16sdp_inst_908.INIT_0 = 16'h0000;
defparam ram16sdp_inst_908.INIT_1 = 16'h0000;
defparam ram16sdp_inst_908.INIT_2 = 16'h0000;
defparam ram16sdp_inst_908.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_909 (
    .DO(ram16sdp_inst_909_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_341),
    .CLK(clk)
);

defparam ram16sdp_inst_909.INIT_0 = 16'h0000;
defparam ram16sdp_inst_909.INIT_1 = 16'h0000;
defparam ram16sdp_inst_909.INIT_2 = 16'h0000;
defparam ram16sdp_inst_909.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_910 (
    .DO(ram16sdp_inst_910_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_341),
    .CLK(clk)
);

defparam ram16sdp_inst_910.INIT_0 = 16'h0000;
defparam ram16sdp_inst_910.INIT_1 = 16'h0000;
defparam ram16sdp_inst_910.INIT_2 = 16'h0000;
defparam ram16sdp_inst_910.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_911 (
    .DO(ram16sdp_inst_911_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_341),
    .CLK(clk)
);

defparam ram16sdp_inst_911.INIT_0 = 16'h0000;
defparam ram16sdp_inst_911.INIT_1 = 16'h0000;
defparam ram16sdp_inst_911.INIT_2 = 16'h0000;
defparam ram16sdp_inst_911.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_912 (
    .DO(ram16sdp_inst_912_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_344),
    .CLK(clk)
);

defparam ram16sdp_inst_912.INIT_0 = 16'h0000;
defparam ram16sdp_inst_912.INIT_1 = 16'h0000;
defparam ram16sdp_inst_912.INIT_2 = 16'h0000;
defparam ram16sdp_inst_912.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_913 (
    .DO(ram16sdp_inst_913_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_344),
    .CLK(clk)
);

defparam ram16sdp_inst_913.INIT_0 = 16'h0000;
defparam ram16sdp_inst_913.INIT_1 = 16'h0000;
defparam ram16sdp_inst_913.INIT_2 = 16'h0000;
defparam ram16sdp_inst_913.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_914 (
    .DO(ram16sdp_inst_914_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_344),
    .CLK(clk)
);

defparam ram16sdp_inst_914.INIT_0 = 16'h0000;
defparam ram16sdp_inst_914.INIT_1 = 16'h0000;
defparam ram16sdp_inst_914.INIT_2 = 16'h0000;
defparam ram16sdp_inst_914.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_915 (
    .DO(ram16sdp_inst_915_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_344),
    .CLK(clk)
);

defparam ram16sdp_inst_915.INIT_0 = 16'h0000;
defparam ram16sdp_inst_915.INIT_1 = 16'h0000;
defparam ram16sdp_inst_915.INIT_2 = 16'h0000;
defparam ram16sdp_inst_915.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_916 (
    .DO(ram16sdp_inst_916_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_344),
    .CLK(clk)
);

defparam ram16sdp_inst_916.INIT_0 = 16'h0000;
defparam ram16sdp_inst_916.INIT_1 = 16'h0000;
defparam ram16sdp_inst_916.INIT_2 = 16'h0000;
defparam ram16sdp_inst_916.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_917 (
    .DO(ram16sdp_inst_917_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_344),
    .CLK(clk)
);

defparam ram16sdp_inst_917.INIT_0 = 16'h0000;
defparam ram16sdp_inst_917.INIT_1 = 16'h0000;
defparam ram16sdp_inst_917.INIT_2 = 16'h0000;
defparam ram16sdp_inst_917.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_918 (
    .DO(ram16sdp_inst_918_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_344),
    .CLK(clk)
);

defparam ram16sdp_inst_918.INIT_0 = 16'h0000;
defparam ram16sdp_inst_918.INIT_1 = 16'h0000;
defparam ram16sdp_inst_918.INIT_2 = 16'h0000;
defparam ram16sdp_inst_918.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_919 (
    .DO(ram16sdp_inst_919_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_344),
    .CLK(clk)
);

defparam ram16sdp_inst_919.INIT_0 = 16'h0000;
defparam ram16sdp_inst_919.INIT_1 = 16'h0000;
defparam ram16sdp_inst_919.INIT_2 = 16'h0000;
defparam ram16sdp_inst_919.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_920 (
    .DO(ram16sdp_inst_920_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16sdp_inst_920.INIT_0 = 16'h0000;
defparam ram16sdp_inst_920.INIT_1 = 16'h0000;
defparam ram16sdp_inst_920.INIT_2 = 16'h0000;
defparam ram16sdp_inst_920.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_921 (
    .DO(ram16sdp_inst_921_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16sdp_inst_921.INIT_0 = 16'h0000;
defparam ram16sdp_inst_921.INIT_1 = 16'h0000;
defparam ram16sdp_inst_921.INIT_2 = 16'h0000;
defparam ram16sdp_inst_921.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_922 (
    .DO(ram16sdp_inst_922_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16sdp_inst_922.INIT_0 = 16'h0000;
defparam ram16sdp_inst_922.INIT_1 = 16'h0000;
defparam ram16sdp_inst_922.INIT_2 = 16'h0000;
defparam ram16sdp_inst_922.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_923 (
    .DO(ram16sdp_inst_923_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16sdp_inst_923.INIT_0 = 16'h0000;
defparam ram16sdp_inst_923.INIT_1 = 16'h0000;
defparam ram16sdp_inst_923.INIT_2 = 16'h0000;
defparam ram16sdp_inst_923.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_924 (
    .DO(ram16sdp_inst_924_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16sdp_inst_924.INIT_0 = 16'h0000;
defparam ram16sdp_inst_924.INIT_1 = 16'h0000;
defparam ram16sdp_inst_924.INIT_2 = 16'h0000;
defparam ram16sdp_inst_924.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_925 (
    .DO(ram16sdp_inst_925_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16sdp_inst_925.INIT_0 = 16'h0000;
defparam ram16sdp_inst_925.INIT_1 = 16'h0000;
defparam ram16sdp_inst_925.INIT_2 = 16'h0000;
defparam ram16sdp_inst_925.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_926 (
    .DO(ram16sdp_inst_926_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16sdp_inst_926.INIT_0 = 16'h0000;
defparam ram16sdp_inst_926.INIT_1 = 16'h0000;
defparam ram16sdp_inst_926.INIT_2 = 16'h0000;
defparam ram16sdp_inst_926.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_927 (
    .DO(ram16sdp_inst_927_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16sdp_inst_927.INIT_0 = 16'h0000;
defparam ram16sdp_inst_927.INIT_1 = 16'h0000;
defparam ram16sdp_inst_927.INIT_2 = 16'h0000;
defparam ram16sdp_inst_927.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_928 (
    .DO(ram16sdp_inst_928_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_350),
    .CLK(clk)
);

defparam ram16sdp_inst_928.INIT_0 = 16'h0000;
defparam ram16sdp_inst_928.INIT_1 = 16'h0000;
defparam ram16sdp_inst_928.INIT_2 = 16'h0000;
defparam ram16sdp_inst_928.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_929 (
    .DO(ram16sdp_inst_929_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_350),
    .CLK(clk)
);

defparam ram16sdp_inst_929.INIT_0 = 16'h0000;
defparam ram16sdp_inst_929.INIT_1 = 16'h0000;
defparam ram16sdp_inst_929.INIT_2 = 16'h0000;
defparam ram16sdp_inst_929.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_930 (
    .DO(ram16sdp_inst_930_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_350),
    .CLK(clk)
);

defparam ram16sdp_inst_930.INIT_0 = 16'h0000;
defparam ram16sdp_inst_930.INIT_1 = 16'h0000;
defparam ram16sdp_inst_930.INIT_2 = 16'h0000;
defparam ram16sdp_inst_930.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_931 (
    .DO(ram16sdp_inst_931_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_350),
    .CLK(clk)
);

defparam ram16sdp_inst_931.INIT_0 = 16'h0000;
defparam ram16sdp_inst_931.INIT_1 = 16'h0000;
defparam ram16sdp_inst_931.INIT_2 = 16'h0000;
defparam ram16sdp_inst_931.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_932 (
    .DO(ram16sdp_inst_932_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_350),
    .CLK(clk)
);

defparam ram16sdp_inst_932.INIT_0 = 16'h0000;
defparam ram16sdp_inst_932.INIT_1 = 16'h0000;
defparam ram16sdp_inst_932.INIT_2 = 16'h0000;
defparam ram16sdp_inst_932.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_933 (
    .DO(ram16sdp_inst_933_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_350),
    .CLK(clk)
);

defparam ram16sdp_inst_933.INIT_0 = 16'h0000;
defparam ram16sdp_inst_933.INIT_1 = 16'h0000;
defparam ram16sdp_inst_933.INIT_2 = 16'h0000;
defparam ram16sdp_inst_933.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_934 (
    .DO(ram16sdp_inst_934_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_350),
    .CLK(clk)
);

defparam ram16sdp_inst_934.INIT_0 = 16'h0000;
defparam ram16sdp_inst_934.INIT_1 = 16'h0000;
defparam ram16sdp_inst_934.INIT_2 = 16'h0000;
defparam ram16sdp_inst_934.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_935 (
    .DO(ram16sdp_inst_935_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_350),
    .CLK(clk)
);

defparam ram16sdp_inst_935.INIT_0 = 16'h0000;
defparam ram16sdp_inst_935.INIT_1 = 16'h0000;
defparam ram16sdp_inst_935.INIT_2 = 16'h0000;
defparam ram16sdp_inst_935.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_936 (
    .DO(ram16sdp_inst_936_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_353),
    .CLK(clk)
);

defparam ram16sdp_inst_936.INIT_0 = 16'h0000;
defparam ram16sdp_inst_936.INIT_1 = 16'h0000;
defparam ram16sdp_inst_936.INIT_2 = 16'h0000;
defparam ram16sdp_inst_936.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_937 (
    .DO(ram16sdp_inst_937_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_353),
    .CLK(clk)
);

defparam ram16sdp_inst_937.INIT_0 = 16'h0000;
defparam ram16sdp_inst_937.INIT_1 = 16'h0000;
defparam ram16sdp_inst_937.INIT_2 = 16'h0000;
defparam ram16sdp_inst_937.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_938 (
    .DO(ram16sdp_inst_938_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_353),
    .CLK(clk)
);

defparam ram16sdp_inst_938.INIT_0 = 16'h0000;
defparam ram16sdp_inst_938.INIT_1 = 16'h0000;
defparam ram16sdp_inst_938.INIT_2 = 16'h0000;
defparam ram16sdp_inst_938.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_939 (
    .DO(ram16sdp_inst_939_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_353),
    .CLK(clk)
);

defparam ram16sdp_inst_939.INIT_0 = 16'h0000;
defparam ram16sdp_inst_939.INIT_1 = 16'h0000;
defparam ram16sdp_inst_939.INIT_2 = 16'h0000;
defparam ram16sdp_inst_939.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_940 (
    .DO(ram16sdp_inst_940_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_353),
    .CLK(clk)
);

defparam ram16sdp_inst_940.INIT_0 = 16'h0000;
defparam ram16sdp_inst_940.INIT_1 = 16'h0000;
defparam ram16sdp_inst_940.INIT_2 = 16'h0000;
defparam ram16sdp_inst_940.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_941 (
    .DO(ram16sdp_inst_941_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_353),
    .CLK(clk)
);

defparam ram16sdp_inst_941.INIT_0 = 16'h0000;
defparam ram16sdp_inst_941.INIT_1 = 16'h0000;
defparam ram16sdp_inst_941.INIT_2 = 16'h0000;
defparam ram16sdp_inst_941.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_942 (
    .DO(ram16sdp_inst_942_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_353),
    .CLK(clk)
);

defparam ram16sdp_inst_942.INIT_0 = 16'h0000;
defparam ram16sdp_inst_942.INIT_1 = 16'h0000;
defparam ram16sdp_inst_942.INIT_2 = 16'h0000;
defparam ram16sdp_inst_942.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_943 (
    .DO(ram16sdp_inst_943_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_353),
    .CLK(clk)
);

defparam ram16sdp_inst_943.INIT_0 = 16'h0000;
defparam ram16sdp_inst_943.INIT_1 = 16'h0000;
defparam ram16sdp_inst_943.INIT_2 = 16'h0000;
defparam ram16sdp_inst_943.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_944 (
    .DO(ram16sdp_inst_944_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_356),
    .CLK(clk)
);

defparam ram16sdp_inst_944.INIT_0 = 16'h0000;
defparam ram16sdp_inst_944.INIT_1 = 16'h0000;
defparam ram16sdp_inst_944.INIT_2 = 16'h0000;
defparam ram16sdp_inst_944.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_945 (
    .DO(ram16sdp_inst_945_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_356),
    .CLK(clk)
);

defparam ram16sdp_inst_945.INIT_0 = 16'h0000;
defparam ram16sdp_inst_945.INIT_1 = 16'h0000;
defparam ram16sdp_inst_945.INIT_2 = 16'h0000;
defparam ram16sdp_inst_945.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_946 (
    .DO(ram16sdp_inst_946_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_356),
    .CLK(clk)
);

defparam ram16sdp_inst_946.INIT_0 = 16'h0000;
defparam ram16sdp_inst_946.INIT_1 = 16'h0000;
defparam ram16sdp_inst_946.INIT_2 = 16'h0000;
defparam ram16sdp_inst_946.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_947 (
    .DO(ram16sdp_inst_947_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_356),
    .CLK(clk)
);

defparam ram16sdp_inst_947.INIT_0 = 16'h0000;
defparam ram16sdp_inst_947.INIT_1 = 16'h0000;
defparam ram16sdp_inst_947.INIT_2 = 16'h0000;
defparam ram16sdp_inst_947.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_948 (
    .DO(ram16sdp_inst_948_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_356),
    .CLK(clk)
);

defparam ram16sdp_inst_948.INIT_0 = 16'h0000;
defparam ram16sdp_inst_948.INIT_1 = 16'h0000;
defparam ram16sdp_inst_948.INIT_2 = 16'h0000;
defparam ram16sdp_inst_948.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_949 (
    .DO(ram16sdp_inst_949_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_356),
    .CLK(clk)
);

defparam ram16sdp_inst_949.INIT_0 = 16'h0000;
defparam ram16sdp_inst_949.INIT_1 = 16'h0000;
defparam ram16sdp_inst_949.INIT_2 = 16'h0000;
defparam ram16sdp_inst_949.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_950 (
    .DO(ram16sdp_inst_950_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_356),
    .CLK(clk)
);

defparam ram16sdp_inst_950.INIT_0 = 16'h0000;
defparam ram16sdp_inst_950.INIT_1 = 16'h0000;
defparam ram16sdp_inst_950.INIT_2 = 16'h0000;
defparam ram16sdp_inst_950.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_951 (
    .DO(ram16sdp_inst_951_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_356),
    .CLK(clk)
);

defparam ram16sdp_inst_951.INIT_0 = 16'h0000;
defparam ram16sdp_inst_951.INIT_1 = 16'h0000;
defparam ram16sdp_inst_951.INIT_2 = 16'h0000;
defparam ram16sdp_inst_951.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_952 (
    .DO(ram16sdp_inst_952_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16sdp_inst_952.INIT_0 = 16'h0000;
defparam ram16sdp_inst_952.INIT_1 = 16'h0000;
defparam ram16sdp_inst_952.INIT_2 = 16'h0000;
defparam ram16sdp_inst_952.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_953 (
    .DO(ram16sdp_inst_953_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16sdp_inst_953.INIT_0 = 16'h0000;
defparam ram16sdp_inst_953.INIT_1 = 16'h0000;
defparam ram16sdp_inst_953.INIT_2 = 16'h0000;
defparam ram16sdp_inst_953.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_954 (
    .DO(ram16sdp_inst_954_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16sdp_inst_954.INIT_0 = 16'h0000;
defparam ram16sdp_inst_954.INIT_1 = 16'h0000;
defparam ram16sdp_inst_954.INIT_2 = 16'h0000;
defparam ram16sdp_inst_954.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_955 (
    .DO(ram16sdp_inst_955_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16sdp_inst_955.INIT_0 = 16'h0000;
defparam ram16sdp_inst_955.INIT_1 = 16'h0000;
defparam ram16sdp_inst_955.INIT_2 = 16'h0000;
defparam ram16sdp_inst_955.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_956 (
    .DO(ram16sdp_inst_956_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16sdp_inst_956.INIT_0 = 16'h0000;
defparam ram16sdp_inst_956.INIT_1 = 16'h0000;
defparam ram16sdp_inst_956.INIT_2 = 16'h0000;
defparam ram16sdp_inst_956.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_957 (
    .DO(ram16sdp_inst_957_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16sdp_inst_957.INIT_0 = 16'h0000;
defparam ram16sdp_inst_957.INIT_1 = 16'h0000;
defparam ram16sdp_inst_957.INIT_2 = 16'h0000;
defparam ram16sdp_inst_957.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_958 (
    .DO(ram16sdp_inst_958_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16sdp_inst_958.INIT_0 = 16'h0000;
defparam ram16sdp_inst_958.INIT_1 = 16'h0000;
defparam ram16sdp_inst_958.INIT_2 = 16'h0000;
defparam ram16sdp_inst_958.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_959 (
    .DO(ram16sdp_inst_959_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16sdp_inst_959.INIT_0 = 16'h0000;
defparam ram16sdp_inst_959.INIT_1 = 16'h0000;
defparam ram16sdp_inst_959.INIT_2 = 16'h0000;
defparam ram16sdp_inst_959.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_960 (
    .DO(ram16sdp_inst_960_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_362),
    .CLK(clk)
);

defparam ram16sdp_inst_960.INIT_0 = 16'h0000;
defparam ram16sdp_inst_960.INIT_1 = 16'h0000;
defparam ram16sdp_inst_960.INIT_2 = 16'h0000;
defparam ram16sdp_inst_960.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_961 (
    .DO(ram16sdp_inst_961_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_362),
    .CLK(clk)
);

defparam ram16sdp_inst_961.INIT_0 = 16'h0000;
defparam ram16sdp_inst_961.INIT_1 = 16'h0000;
defparam ram16sdp_inst_961.INIT_2 = 16'h0000;
defparam ram16sdp_inst_961.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_962 (
    .DO(ram16sdp_inst_962_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_362),
    .CLK(clk)
);

defparam ram16sdp_inst_962.INIT_0 = 16'h0000;
defparam ram16sdp_inst_962.INIT_1 = 16'h0000;
defparam ram16sdp_inst_962.INIT_2 = 16'h0000;
defparam ram16sdp_inst_962.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_963 (
    .DO(ram16sdp_inst_963_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_362),
    .CLK(clk)
);

defparam ram16sdp_inst_963.INIT_0 = 16'h0000;
defparam ram16sdp_inst_963.INIT_1 = 16'h0000;
defparam ram16sdp_inst_963.INIT_2 = 16'h0000;
defparam ram16sdp_inst_963.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_964 (
    .DO(ram16sdp_inst_964_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_362),
    .CLK(clk)
);

defparam ram16sdp_inst_964.INIT_0 = 16'h0000;
defparam ram16sdp_inst_964.INIT_1 = 16'h0000;
defparam ram16sdp_inst_964.INIT_2 = 16'h0000;
defparam ram16sdp_inst_964.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_965 (
    .DO(ram16sdp_inst_965_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_362),
    .CLK(clk)
);

defparam ram16sdp_inst_965.INIT_0 = 16'h0000;
defparam ram16sdp_inst_965.INIT_1 = 16'h0000;
defparam ram16sdp_inst_965.INIT_2 = 16'h0000;
defparam ram16sdp_inst_965.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_966 (
    .DO(ram16sdp_inst_966_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_362),
    .CLK(clk)
);

defparam ram16sdp_inst_966.INIT_0 = 16'h0000;
defparam ram16sdp_inst_966.INIT_1 = 16'h0000;
defparam ram16sdp_inst_966.INIT_2 = 16'h0000;
defparam ram16sdp_inst_966.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_967 (
    .DO(ram16sdp_inst_967_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_362),
    .CLK(clk)
);

defparam ram16sdp_inst_967.INIT_0 = 16'h0000;
defparam ram16sdp_inst_967.INIT_1 = 16'h0000;
defparam ram16sdp_inst_967.INIT_2 = 16'h0000;
defparam ram16sdp_inst_967.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_968 (
    .DO(ram16sdp_inst_968_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_365),
    .CLK(clk)
);

defparam ram16sdp_inst_968.INIT_0 = 16'h0000;
defparam ram16sdp_inst_968.INIT_1 = 16'h0000;
defparam ram16sdp_inst_968.INIT_2 = 16'h0000;
defparam ram16sdp_inst_968.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_969 (
    .DO(ram16sdp_inst_969_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_365),
    .CLK(clk)
);

defparam ram16sdp_inst_969.INIT_0 = 16'h0000;
defparam ram16sdp_inst_969.INIT_1 = 16'h0000;
defparam ram16sdp_inst_969.INIT_2 = 16'h0000;
defparam ram16sdp_inst_969.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_970 (
    .DO(ram16sdp_inst_970_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_365),
    .CLK(clk)
);

defparam ram16sdp_inst_970.INIT_0 = 16'h0000;
defparam ram16sdp_inst_970.INIT_1 = 16'h0000;
defparam ram16sdp_inst_970.INIT_2 = 16'h0000;
defparam ram16sdp_inst_970.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_971 (
    .DO(ram16sdp_inst_971_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_365),
    .CLK(clk)
);

defparam ram16sdp_inst_971.INIT_0 = 16'h0000;
defparam ram16sdp_inst_971.INIT_1 = 16'h0000;
defparam ram16sdp_inst_971.INIT_2 = 16'h0000;
defparam ram16sdp_inst_971.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_972 (
    .DO(ram16sdp_inst_972_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_365),
    .CLK(clk)
);

defparam ram16sdp_inst_972.INIT_0 = 16'h0000;
defparam ram16sdp_inst_972.INIT_1 = 16'h0000;
defparam ram16sdp_inst_972.INIT_2 = 16'h0000;
defparam ram16sdp_inst_972.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_973 (
    .DO(ram16sdp_inst_973_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_365),
    .CLK(clk)
);

defparam ram16sdp_inst_973.INIT_0 = 16'h0000;
defparam ram16sdp_inst_973.INIT_1 = 16'h0000;
defparam ram16sdp_inst_973.INIT_2 = 16'h0000;
defparam ram16sdp_inst_973.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_974 (
    .DO(ram16sdp_inst_974_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_365),
    .CLK(clk)
);

defparam ram16sdp_inst_974.INIT_0 = 16'h0000;
defparam ram16sdp_inst_974.INIT_1 = 16'h0000;
defparam ram16sdp_inst_974.INIT_2 = 16'h0000;
defparam ram16sdp_inst_974.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_975 (
    .DO(ram16sdp_inst_975_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_365),
    .CLK(clk)
);

defparam ram16sdp_inst_975.INIT_0 = 16'h0000;
defparam ram16sdp_inst_975.INIT_1 = 16'h0000;
defparam ram16sdp_inst_975.INIT_2 = 16'h0000;
defparam ram16sdp_inst_975.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_976 (
    .DO(ram16sdp_inst_976_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_368),
    .CLK(clk)
);

defparam ram16sdp_inst_976.INIT_0 = 16'h0000;
defparam ram16sdp_inst_976.INIT_1 = 16'h0000;
defparam ram16sdp_inst_976.INIT_2 = 16'h0000;
defparam ram16sdp_inst_976.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_977 (
    .DO(ram16sdp_inst_977_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_368),
    .CLK(clk)
);

defparam ram16sdp_inst_977.INIT_0 = 16'h0000;
defparam ram16sdp_inst_977.INIT_1 = 16'h0000;
defparam ram16sdp_inst_977.INIT_2 = 16'h0000;
defparam ram16sdp_inst_977.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_978 (
    .DO(ram16sdp_inst_978_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_368),
    .CLK(clk)
);

defparam ram16sdp_inst_978.INIT_0 = 16'h0000;
defparam ram16sdp_inst_978.INIT_1 = 16'h0000;
defparam ram16sdp_inst_978.INIT_2 = 16'h0000;
defparam ram16sdp_inst_978.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_979 (
    .DO(ram16sdp_inst_979_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_368),
    .CLK(clk)
);

defparam ram16sdp_inst_979.INIT_0 = 16'h0000;
defparam ram16sdp_inst_979.INIT_1 = 16'h0000;
defparam ram16sdp_inst_979.INIT_2 = 16'h0000;
defparam ram16sdp_inst_979.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_980 (
    .DO(ram16sdp_inst_980_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_368),
    .CLK(clk)
);

defparam ram16sdp_inst_980.INIT_0 = 16'h0000;
defparam ram16sdp_inst_980.INIT_1 = 16'h0000;
defparam ram16sdp_inst_980.INIT_2 = 16'h0000;
defparam ram16sdp_inst_980.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_981 (
    .DO(ram16sdp_inst_981_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_368),
    .CLK(clk)
);

defparam ram16sdp_inst_981.INIT_0 = 16'h0000;
defparam ram16sdp_inst_981.INIT_1 = 16'h0000;
defparam ram16sdp_inst_981.INIT_2 = 16'h0000;
defparam ram16sdp_inst_981.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_982 (
    .DO(ram16sdp_inst_982_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_368),
    .CLK(clk)
);

defparam ram16sdp_inst_982.INIT_0 = 16'h0000;
defparam ram16sdp_inst_982.INIT_1 = 16'h0000;
defparam ram16sdp_inst_982.INIT_2 = 16'h0000;
defparam ram16sdp_inst_982.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_983 (
    .DO(ram16sdp_inst_983_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_368),
    .CLK(clk)
);

defparam ram16sdp_inst_983.INIT_0 = 16'h0000;
defparam ram16sdp_inst_983.INIT_1 = 16'h0000;
defparam ram16sdp_inst_983.INIT_2 = 16'h0000;
defparam ram16sdp_inst_983.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_984 (
    .DO(ram16sdp_inst_984_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16sdp_inst_984.INIT_0 = 16'h0000;
defparam ram16sdp_inst_984.INIT_1 = 16'h0000;
defparam ram16sdp_inst_984.INIT_2 = 16'h0000;
defparam ram16sdp_inst_984.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_985 (
    .DO(ram16sdp_inst_985_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16sdp_inst_985.INIT_0 = 16'h0000;
defparam ram16sdp_inst_985.INIT_1 = 16'h0000;
defparam ram16sdp_inst_985.INIT_2 = 16'h0000;
defparam ram16sdp_inst_985.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_986 (
    .DO(ram16sdp_inst_986_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16sdp_inst_986.INIT_0 = 16'h0000;
defparam ram16sdp_inst_986.INIT_1 = 16'h0000;
defparam ram16sdp_inst_986.INIT_2 = 16'h0000;
defparam ram16sdp_inst_986.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_987 (
    .DO(ram16sdp_inst_987_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16sdp_inst_987.INIT_0 = 16'h0000;
defparam ram16sdp_inst_987.INIT_1 = 16'h0000;
defparam ram16sdp_inst_987.INIT_2 = 16'h0000;
defparam ram16sdp_inst_987.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_988 (
    .DO(ram16sdp_inst_988_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16sdp_inst_988.INIT_0 = 16'h0000;
defparam ram16sdp_inst_988.INIT_1 = 16'h0000;
defparam ram16sdp_inst_988.INIT_2 = 16'h0000;
defparam ram16sdp_inst_988.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_989 (
    .DO(ram16sdp_inst_989_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16sdp_inst_989.INIT_0 = 16'h0000;
defparam ram16sdp_inst_989.INIT_1 = 16'h0000;
defparam ram16sdp_inst_989.INIT_2 = 16'h0000;
defparam ram16sdp_inst_989.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_990 (
    .DO(ram16sdp_inst_990_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16sdp_inst_990.INIT_0 = 16'h0000;
defparam ram16sdp_inst_990.INIT_1 = 16'h0000;
defparam ram16sdp_inst_990.INIT_2 = 16'h0000;
defparam ram16sdp_inst_990.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_991 (
    .DO(ram16sdp_inst_991_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16sdp_inst_991.INIT_0 = 16'h0000;
defparam ram16sdp_inst_991.INIT_1 = 16'h0000;
defparam ram16sdp_inst_991.INIT_2 = 16'h0000;
defparam ram16sdp_inst_991.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_992 (
    .DO(ram16sdp_inst_992_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_374),
    .CLK(clk)
);

defparam ram16sdp_inst_992.INIT_0 = 16'h0000;
defparam ram16sdp_inst_992.INIT_1 = 16'h0000;
defparam ram16sdp_inst_992.INIT_2 = 16'h0000;
defparam ram16sdp_inst_992.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_993 (
    .DO(ram16sdp_inst_993_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_374),
    .CLK(clk)
);

defparam ram16sdp_inst_993.INIT_0 = 16'h0000;
defparam ram16sdp_inst_993.INIT_1 = 16'h0000;
defparam ram16sdp_inst_993.INIT_2 = 16'h0000;
defparam ram16sdp_inst_993.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_994 (
    .DO(ram16sdp_inst_994_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_374),
    .CLK(clk)
);

defparam ram16sdp_inst_994.INIT_0 = 16'h0000;
defparam ram16sdp_inst_994.INIT_1 = 16'h0000;
defparam ram16sdp_inst_994.INIT_2 = 16'h0000;
defparam ram16sdp_inst_994.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_995 (
    .DO(ram16sdp_inst_995_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_374),
    .CLK(clk)
);

defparam ram16sdp_inst_995.INIT_0 = 16'h0000;
defparam ram16sdp_inst_995.INIT_1 = 16'h0000;
defparam ram16sdp_inst_995.INIT_2 = 16'h0000;
defparam ram16sdp_inst_995.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_996 (
    .DO(ram16sdp_inst_996_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_374),
    .CLK(clk)
);

defparam ram16sdp_inst_996.INIT_0 = 16'h0000;
defparam ram16sdp_inst_996.INIT_1 = 16'h0000;
defparam ram16sdp_inst_996.INIT_2 = 16'h0000;
defparam ram16sdp_inst_996.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_997 (
    .DO(ram16sdp_inst_997_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_374),
    .CLK(clk)
);

defparam ram16sdp_inst_997.INIT_0 = 16'h0000;
defparam ram16sdp_inst_997.INIT_1 = 16'h0000;
defparam ram16sdp_inst_997.INIT_2 = 16'h0000;
defparam ram16sdp_inst_997.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_998 (
    .DO(ram16sdp_inst_998_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_374),
    .CLK(clk)
);

defparam ram16sdp_inst_998.INIT_0 = 16'h0000;
defparam ram16sdp_inst_998.INIT_1 = 16'h0000;
defparam ram16sdp_inst_998.INIT_2 = 16'h0000;
defparam ram16sdp_inst_998.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_999 (
    .DO(ram16sdp_inst_999_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_374),
    .CLK(clk)
);

defparam ram16sdp_inst_999.INIT_0 = 16'h0000;
defparam ram16sdp_inst_999.INIT_1 = 16'h0000;
defparam ram16sdp_inst_999.INIT_2 = 16'h0000;
defparam ram16sdp_inst_999.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1000 (
    .DO(ram16sdp_inst_1000_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_377),
    .CLK(clk)
);

defparam ram16sdp_inst_1000.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1000.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1000.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1000.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1001 (
    .DO(ram16sdp_inst_1001_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_377),
    .CLK(clk)
);

defparam ram16sdp_inst_1001.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1001.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1001.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1001.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1002 (
    .DO(ram16sdp_inst_1002_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_377),
    .CLK(clk)
);

defparam ram16sdp_inst_1002.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1002.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1002.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1002.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1003 (
    .DO(ram16sdp_inst_1003_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_377),
    .CLK(clk)
);

defparam ram16sdp_inst_1003.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1003.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1003.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1003.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1004 (
    .DO(ram16sdp_inst_1004_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_377),
    .CLK(clk)
);

defparam ram16sdp_inst_1004.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1004.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1004.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1004.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1005 (
    .DO(ram16sdp_inst_1005_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_377),
    .CLK(clk)
);

defparam ram16sdp_inst_1005.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1005.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1005.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1005.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1006 (
    .DO(ram16sdp_inst_1006_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_377),
    .CLK(clk)
);

defparam ram16sdp_inst_1006.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1006.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1006.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1006.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1007 (
    .DO(ram16sdp_inst_1007_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_377),
    .CLK(clk)
);

defparam ram16sdp_inst_1007.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1007.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1007.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1007.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1008 (
    .DO(ram16sdp_inst_1008_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_380),
    .CLK(clk)
);

defparam ram16sdp_inst_1008.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1008.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1008.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1008.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1009 (
    .DO(ram16sdp_inst_1009_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_380),
    .CLK(clk)
);

defparam ram16sdp_inst_1009.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1009.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1009.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1009.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1010 (
    .DO(ram16sdp_inst_1010_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_380),
    .CLK(clk)
);

defparam ram16sdp_inst_1010.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1010.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1010.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1010.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1011 (
    .DO(ram16sdp_inst_1011_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_380),
    .CLK(clk)
);

defparam ram16sdp_inst_1011.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1011.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1011.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1011.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1012 (
    .DO(ram16sdp_inst_1012_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_380),
    .CLK(clk)
);

defparam ram16sdp_inst_1012.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1012.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1012.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1012.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1013 (
    .DO(ram16sdp_inst_1013_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_380),
    .CLK(clk)
);

defparam ram16sdp_inst_1013.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1013.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1013.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1013.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1014 (
    .DO(ram16sdp_inst_1014_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_380),
    .CLK(clk)
);

defparam ram16sdp_inst_1014.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1014.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1014.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1014.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1015 (
    .DO(ram16sdp_inst_1015_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_380),
    .CLK(clk)
);

defparam ram16sdp_inst_1015.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1015.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1015.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1015.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1016 (
    .DO(ram16sdp_inst_1016_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16sdp_inst_1016.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1016.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1016.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1016.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1017 (
    .DO(ram16sdp_inst_1017_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16sdp_inst_1017.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1017.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1017.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1017.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1018 (
    .DO(ram16sdp_inst_1018_dout[11:8]),
    .DI(di[11:8]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16sdp_inst_1018.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1018.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1018.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1018.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1019 (
    .DO(ram16sdp_inst_1019_dout[15:12]),
    .DI(di[15:12]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16sdp_inst_1019.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1019.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1019.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1019.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1020 (
    .DO(ram16sdp_inst_1020_dout[19:16]),
    .DI(di[19:16]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16sdp_inst_1020.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1020.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1020.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1020.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1021 (
    .DO(ram16sdp_inst_1021_dout[23:20]),
    .DI(di[23:20]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16sdp_inst_1021.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1021.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1021.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1021.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1022 (
    .DO(ram16sdp_inst_1022_dout[27:24]),
    .DI(di[27:24]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16sdp_inst_1022.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1022.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1022.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1022.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1023 (
    .DO(ram16sdp_inst_1023_dout[31:28]),
    .DI(di[31:28]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16sdp_inst_1023.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1023.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1023.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1023.INIT_3 = 16'h0000;

MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(ram16sdp_inst_0_dout[0]),
  .I1(ram16sdp_inst_8_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(ram16sdp_inst_16_dout[0]),
  .I1(ram16sdp_inst_24_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(ram16sdp_inst_32_dout[0]),
  .I1(ram16sdp_inst_40_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(ram16sdp_inst_48_dout[0]),
  .I1(ram16sdp_inst_56_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(ram16sdp_inst_64_dout[0]),
  .I1(ram16sdp_inst_72_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(ram16sdp_inst_80_dout[0]),
  .I1(ram16sdp_inst_88_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(ram16sdp_inst_96_dout[0]),
  .I1(ram16sdp_inst_104_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(ram16sdp_inst_112_dout[0]),
  .I1(ram16sdp_inst_120_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(ram16sdp_inst_128_dout[0]),
  .I1(ram16sdp_inst_136_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(ram16sdp_inst_144_dout[0]),
  .I1(ram16sdp_inst_152_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(ram16sdp_inst_160_dout[0]),
  .I1(ram16sdp_inst_168_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(ram16sdp_inst_176_dout[0]),
  .I1(ram16sdp_inst_184_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(ram16sdp_inst_192_dout[0]),
  .I1(ram16sdp_inst_200_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(ram16sdp_inst_208_dout[0]),
  .I1(ram16sdp_inst_216_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(ram16sdp_inst_224_dout[0]),
  .I1(ram16sdp_inst_232_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(ram16sdp_inst_240_dout[0]),
  .I1(ram16sdp_inst_248_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(ram16sdp_inst_256_dout[0]),
  .I1(ram16sdp_inst_264_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(ram16sdp_inst_272_dout[0]),
  .I1(ram16sdp_inst_280_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(ram16sdp_inst_288_dout[0]),
  .I1(ram16sdp_inst_296_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(ram16sdp_inst_304_dout[0]),
  .I1(ram16sdp_inst_312_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(ram16sdp_inst_320_dout[0]),
  .I1(ram16sdp_inst_328_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(ram16sdp_inst_336_dout[0]),
  .I1(ram16sdp_inst_344_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(ram16sdp_inst_352_dout[0]),
  .I1(ram16sdp_inst_360_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(ram16sdp_inst_368_dout[0]),
  .I1(ram16sdp_inst_376_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(ram16sdp_inst_384_dout[0]),
  .I1(ram16sdp_inst_392_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(ram16sdp_inst_400_dout[0]),
  .I1(ram16sdp_inst_408_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(ram16sdp_inst_416_dout[0]),
  .I1(ram16sdp_inst_424_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(ram16sdp_inst_432_dout[0]),
  .I1(ram16sdp_inst_440_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(ram16sdp_inst_448_dout[0]),
  .I1(ram16sdp_inst_456_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(ram16sdp_inst_464_dout[0]),
  .I1(ram16sdp_inst_472_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(ram16sdp_inst_480_dout[0]),
  .I1(ram16sdp_inst_488_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(ram16sdp_inst_496_dout[0]),
  .I1(ram16sdp_inst_504_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(ram16sdp_inst_512_dout[0]),
  .I1(ram16sdp_inst_520_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(ram16sdp_inst_528_dout[0]),
  .I1(ram16sdp_inst_536_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(ram16sdp_inst_544_dout[0]),
  .I1(ram16sdp_inst_552_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(ram16sdp_inst_560_dout[0]),
  .I1(ram16sdp_inst_568_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(ram16sdp_inst_576_dout[0]),
  .I1(ram16sdp_inst_584_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(ram16sdp_inst_592_dout[0]),
  .I1(ram16sdp_inst_600_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(ram16sdp_inst_608_dout[0]),
  .I1(ram16sdp_inst_616_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(ram16sdp_inst_624_dout[0]),
  .I1(ram16sdp_inst_632_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(ram16sdp_inst_640_dout[0]),
  .I1(ram16sdp_inst_648_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(ram16sdp_inst_656_dout[0]),
  .I1(ram16sdp_inst_664_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(ram16sdp_inst_672_dout[0]),
  .I1(ram16sdp_inst_680_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(ram16sdp_inst_688_dout[0]),
  .I1(ram16sdp_inst_696_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(ram16sdp_inst_704_dout[0]),
  .I1(ram16sdp_inst_712_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(ram16sdp_inst_720_dout[0]),
  .I1(ram16sdp_inst_728_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(ram16sdp_inst_736_dout[0]),
  .I1(ram16sdp_inst_744_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(ram16sdp_inst_752_dout[0]),
  .I1(ram16sdp_inst_760_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(ram16sdp_inst_768_dout[0]),
  .I1(ram16sdp_inst_776_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(ram16sdp_inst_784_dout[0]),
  .I1(ram16sdp_inst_792_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(ram16sdp_inst_800_dout[0]),
  .I1(ram16sdp_inst_808_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(ram16sdp_inst_816_dout[0]),
  .I1(ram16sdp_inst_824_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(ram16sdp_inst_832_dout[0]),
  .I1(ram16sdp_inst_840_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(ram16sdp_inst_848_dout[0]),
  .I1(ram16sdp_inst_856_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(ram16sdp_inst_864_dout[0]),
  .I1(ram16sdp_inst_872_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(ram16sdp_inst_880_dout[0]),
  .I1(ram16sdp_inst_888_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(ram16sdp_inst_896_dout[0]),
  .I1(ram16sdp_inst_904_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(ram16sdp_inst_912_dout[0]),
  .I1(ram16sdp_inst_920_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(ram16sdp_inst_928_dout[0]),
  .I1(ram16sdp_inst_936_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(ram16sdp_inst_944_dout[0]),
  .I1(ram16sdp_inst_952_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(ram16sdp_inst_960_dout[0]),
  .I1(ram16sdp_inst_968_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(ram16sdp_inst_976_dout[0]),
  .I1(ram16sdp_inst_984_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(ram16sdp_inst_992_dout[0]),
  .I1(ram16sdp_inst_1000_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(ram16sdp_inst_1008_dout[0]),
  .I1(ram16sdp_inst_1016_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(rad[5])
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(rad[5])
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(rad[5])
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(rad[5])
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(rad[5])
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(rad[5])
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(rad[5])
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(rad[5])
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(rad[5])
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(rad[5])
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(rad[5])
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(rad[5])
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(rad[5])
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(rad[5])
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(rad[5])
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(rad[5])
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(rad[5])
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(rad[5])
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(rad[5])
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(rad[5])
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(rad[5])
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(rad[5])
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_44),
  .I1(mux_o_45),
  .S0(rad[5])
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_46),
  .I1(mux_o_47),
  .S0(rad[5])
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_48),
  .I1(mux_o_49),
  .S0(rad[5])
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_50),
  .I1(mux_o_51),
  .S0(rad[5])
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_52),
  .I1(mux_o_53),
  .S0(rad[5])
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_54),
  .I1(mux_o_55),
  .S0(rad[5])
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(rad[5])
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(rad[5])
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(rad[5])
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(rad[5])
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(rad[6])
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(rad[6])
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(rad[6])
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(rad[6])
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(rad[6])
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(rad[6])
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_76),
  .I1(mux_o_77),
  .S0(rad[6])
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_78),
  .I1(mux_o_79),
  .S0(rad[6])
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(mux_o_80),
  .I1(mux_o_81),
  .S0(rad[6])
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(mux_o_82),
  .I1(mux_o_83),
  .S0(rad[6])
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(rad[6])
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(rad[6])
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(rad[6])
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(rad[6])
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(rad[6])
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(rad[6])
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(rad[7])
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(rad[7])
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(rad[7])
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(rad[7])
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_104),
  .I1(mux_o_105),
  .S0(rad[7])
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_106),
  .I1(mux_o_107),
  .S0(rad[7])
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_108),
  .I1(mux_o_109),
  .S0(rad[7])
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_110),
  .I1(mux_o_111),
  .S0(rad[7])
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(rad[8])
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_114),
  .I1(mux_o_115),
  .S0(rad[8])
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(mux_o_116),
  .I1(mux_o_117),
  .S0(rad[8])
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(mux_o_118),
  .I1(mux_o_119),
  .S0(rad[8])
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(mux_o_120),
  .I1(mux_o_121),
  .S0(rad[9])
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(mux_o_122),
  .I1(mux_o_123),
  .S0(rad[9])
);
MUX2 mux_inst_126 (
  .O(dout[0]),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(rad[10])
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(ram16sdp_inst_0_dout[1]),
  .I1(ram16sdp_inst_8_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(ram16sdp_inst_16_dout[1]),
  .I1(ram16sdp_inst_24_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(ram16sdp_inst_32_dout[1]),
  .I1(ram16sdp_inst_40_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(ram16sdp_inst_48_dout[1]),
  .I1(ram16sdp_inst_56_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(ram16sdp_inst_64_dout[1]),
  .I1(ram16sdp_inst_72_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(ram16sdp_inst_80_dout[1]),
  .I1(ram16sdp_inst_88_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(ram16sdp_inst_96_dout[1]),
  .I1(ram16sdp_inst_104_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(ram16sdp_inst_112_dout[1]),
  .I1(ram16sdp_inst_120_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(ram16sdp_inst_128_dout[1]),
  .I1(ram16sdp_inst_136_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(ram16sdp_inst_144_dout[1]),
  .I1(ram16sdp_inst_152_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(ram16sdp_inst_160_dout[1]),
  .I1(ram16sdp_inst_168_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(ram16sdp_inst_176_dout[1]),
  .I1(ram16sdp_inst_184_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(ram16sdp_inst_192_dout[1]),
  .I1(ram16sdp_inst_200_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(ram16sdp_inst_208_dout[1]),
  .I1(ram16sdp_inst_216_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(ram16sdp_inst_224_dout[1]),
  .I1(ram16sdp_inst_232_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(ram16sdp_inst_240_dout[1]),
  .I1(ram16sdp_inst_248_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(ram16sdp_inst_256_dout[1]),
  .I1(ram16sdp_inst_264_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(ram16sdp_inst_272_dout[1]),
  .I1(ram16sdp_inst_280_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(ram16sdp_inst_288_dout[1]),
  .I1(ram16sdp_inst_296_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(ram16sdp_inst_304_dout[1]),
  .I1(ram16sdp_inst_312_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(ram16sdp_inst_320_dout[1]),
  .I1(ram16sdp_inst_328_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(ram16sdp_inst_336_dout[1]),
  .I1(ram16sdp_inst_344_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(ram16sdp_inst_352_dout[1]),
  .I1(ram16sdp_inst_360_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(ram16sdp_inst_368_dout[1]),
  .I1(ram16sdp_inst_376_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(ram16sdp_inst_384_dout[1]),
  .I1(ram16sdp_inst_392_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(ram16sdp_inst_400_dout[1]),
  .I1(ram16sdp_inst_408_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(ram16sdp_inst_416_dout[1]),
  .I1(ram16sdp_inst_424_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(ram16sdp_inst_432_dout[1]),
  .I1(ram16sdp_inst_440_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(ram16sdp_inst_448_dout[1]),
  .I1(ram16sdp_inst_456_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(ram16sdp_inst_464_dout[1]),
  .I1(ram16sdp_inst_472_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(ram16sdp_inst_480_dout[1]),
  .I1(ram16sdp_inst_488_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(ram16sdp_inst_496_dout[1]),
  .I1(ram16sdp_inst_504_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(ram16sdp_inst_512_dout[1]),
  .I1(ram16sdp_inst_520_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(ram16sdp_inst_528_dout[1]),
  .I1(ram16sdp_inst_536_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(ram16sdp_inst_544_dout[1]),
  .I1(ram16sdp_inst_552_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(ram16sdp_inst_560_dout[1]),
  .I1(ram16sdp_inst_568_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(ram16sdp_inst_576_dout[1]),
  .I1(ram16sdp_inst_584_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(ram16sdp_inst_592_dout[1]),
  .I1(ram16sdp_inst_600_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(ram16sdp_inst_608_dout[1]),
  .I1(ram16sdp_inst_616_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(ram16sdp_inst_624_dout[1]),
  .I1(ram16sdp_inst_632_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(ram16sdp_inst_640_dout[1]),
  .I1(ram16sdp_inst_648_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(ram16sdp_inst_656_dout[1]),
  .I1(ram16sdp_inst_664_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(ram16sdp_inst_672_dout[1]),
  .I1(ram16sdp_inst_680_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(ram16sdp_inst_688_dout[1]),
  .I1(ram16sdp_inst_696_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(ram16sdp_inst_704_dout[1]),
  .I1(ram16sdp_inst_712_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(ram16sdp_inst_720_dout[1]),
  .I1(ram16sdp_inst_728_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(ram16sdp_inst_736_dout[1]),
  .I1(ram16sdp_inst_744_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(ram16sdp_inst_752_dout[1]),
  .I1(ram16sdp_inst_760_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(ram16sdp_inst_768_dout[1]),
  .I1(ram16sdp_inst_776_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(ram16sdp_inst_784_dout[1]),
  .I1(ram16sdp_inst_792_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(ram16sdp_inst_800_dout[1]),
  .I1(ram16sdp_inst_808_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(ram16sdp_inst_816_dout[1]),
  .I1(ram16sdp_inst_824_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(ram16sdp_inst_832_dout[1]),
  .I1(ram16sdp_inst_840_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(ram16sdp_inst_848_dout[1]),
  .I1(ram16sdp_inst_856_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(ram16sdp_inst_864_dout[1]),
  .I1(ram16sdp_inst_872_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(ram16sdp_inst_880_dout[1]),
  .I1(ram16sdp_inst_888_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(ram16sdp_inst_896_dout[1]),
  .I1(ram16sdp_inst_904_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(ram16sdp_inst_912_dout[1]),
  .I1(ram16sdp_inst_920_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(ram16sdp_inst_928_dout[1]),
  .I1(ram16sdp_inst_936_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(ram16sdp_inst_944_dout[1]),
  .I1(ram16sdp_inst_952_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(ram16sdp_inst_960_dout[1]),
  .I1(ram16sdp_inst_968_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(ram16sdp_inst_976_dout[1]),
  .I1(ram16sdp_inst_984_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(ram16sdp_inst_992_dout[1]),
  .I1(ram16sdp_inst_1000_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(ram16sdp_inst_1008_dout[1]),
  .I1(ram16sdp_inst_1016_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(mux_o_127),
  .I1(mux_o_128),
  .S0(rad[5])
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(mux_o_129),
  .I1(mux_o_130),
  .S0(rad[5])
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_131),
  .I1(mux_o_132),
  .S0(rad[5])
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(rad[5])
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(rad[5])
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(rad[5])
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(rad[5])
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(mux_o_141),
  .I1(mux_o_142),
  .S0(rad[5])
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(mux_o_143),
  .I1(mux_o_144),
  .S0(rad[5])
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(mux_o_145),
  .I1(mux_o_146),
  .S0(rad[5])
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(rad[5])
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(mux_o_149),
  .I1(mux_o_150),
  .S0(rad[5])
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_151),
  .I1(mux_o_152),
  .S0(rad[5])
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_153),
  .I1(mux_o_154),
  .S0(rad[5])
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_155),
  .I1(mux_o_156),
  .S0(rad[5])
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_157),
  .I1(mux_o_158),
  .S0(rad[5])
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_159),
  .I1(mux_o_160),
  .S0(rad[5])
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(rad[5])
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(mux_o_163),
  .I1(mux_o_164),
  .S0(rad[5])
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(rad[5])
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(rad[5])
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(rad[5])
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(rad[5])
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(rad[5])
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(rad[5])
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(rad[5])
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(rad[5])
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(rad[5])
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(rad[5])
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(mux_o_185),
  .I1(mux_o_186),
  .S0(rad[5])
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_187),
  .I1(mux_o_188),
  .S0(rad[5])
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(rad[5])
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(rad[6])
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(mux_o_193),
  .I1(mux_o_194),
  .S0(rad[6])
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(mux_o_195),
  .I1(mux_o_196),
  .S0(rad[6])
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(mux_o_197),
  .I1(mux_o_198),
  .S0(rad[6])
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(mux_o_199),
  .I1(mux_o_200),
  .S0(rad[6])
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(rad[6])
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(rad[6])
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(rad[6])
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(rad[6])
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(mux_o_209),
  .I1(mux_o_210),
  .S0(rad[6])
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_211),
  .I1(mux_o_212),
  .S0(rad[6])
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_213),
  .I1(mux_o_214),
  .S0(rad[6])
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_215),
  .I1(mux_o_216),
  .S0(rad[6])
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(rad[6])
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(rad[6])
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(rad[6])
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_223),
  .I1(mux_o_224),
  .S0(rad[7])
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(rad[7])
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(rad[7])
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(rad[7])
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(rad[7])
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(rad[7])
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(rad[7])
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(rad[7])
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(rad[8])
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(rad[8])
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(rad[8])
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(rad[8])
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(mux_o_247),
  .I1(mux_o_248),
  .S0(rad[9])
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(mux_o_249),
  .I1(mux_o_250),
  .S0(rad[9])
);
MUX2 mux_inst_253 (
  .O(dout[1]),
  .I0(mux_o_251),
  .I1(mux_o_252),
  .S0(rad[10])
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(ram16sdp_inst_0_dout[2]),
  .I1(ram16sdp_inst_8_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(ram16sdp_inst_16_dout[2]),
  .I1(ram16sdp_inst_24_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(ram16sdp_inst_32_dout[2]),
  .I1(ram16sdp_inst_40_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(ram16sdp_inst_48_dout[2]),
  .I1(ram16sdp_inst_56_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(ram16sdp_inst_64_dout[2]),
  .I1(ram16sdp_inst_72_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(ram16sdp_inst_80_dout[2]),
  .I1(ram16sdp_inst_88_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(ram16sdp_inst_96_dout[2]),
  .I1(ram16sdp_inst_104_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(ram16sdp_inst_112_dout[2]),
  .I1(ram16sdp_inst_120_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(ram16sdp_inst_128_dout[2]),
  .I1(ram16sdp_inst_136_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(ram16sdp_inst_144_dout[2]),
  .I1(ram16sdp_inst_152_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(ram16sdp_inst_160_dout[2]),
  .I1(ram16sdp_inst_168_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(ram16sdp_inst_176_dout[2]),
  .I1(ram16sdp_inst_184_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(ram16sdp_inst_192_dout[2]),
  .I1(ram16sdp_inst_200_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(ram16sdp_inst_208_dout[2]),
  .I1(ram16sdp_inst_216_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(ram16sdp_inst_224_dout[2]),
  .I1(ram16sdp_inst_232_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(ram16sdp_inst_240_dout[2]),
  .I1(ram16sdp_inst_248_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(ram16sdp_inst_256_dout[2]),
  .I1(ram16sdp_inst_264_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(ram16sdp_inst_272_dout[2]),
  .I1(ram16sdp_inst_280_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(ram16sdp_inst_288_dout[2]),
  .I1(ram16sdp_inst_296_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(ram16sdp_inst_304_dout[2]),
  .I1(ram16sdp_inst_312_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(ram16sdp_inst_320_dout[2]),
  .I1(ram16sdp_inst_328_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(ram16sdp_inst_336_dout[2]),
  .I1(ram16sdp_inst_344_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(ram16sdp_inst_352_dout[2]),
  .I1(ram16sdp_inst_360_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(ram16sdp_inst_368_dout[2]),
  .I1(ram16sdp_inst_376_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(ram16sdp_inst_384_dout[2]),
  .I1(ram16sdp_inst_392_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(ram16sdp_inst_400_dout[2]),
  .I1(ram16sdp_inst_408_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(ram16sdp_inst_416_dout[2]),
  .I1(ram16sdp_inst_424_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(ram16sdp_inst_432_dout[2]),
  .I1(ram16sdp_inst_440_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(ram16sdp_inst_448_dout[2]),
  .I1(ram16sdp_inst_456_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(ram16sdp_inst_464_dout[2]),
  .I1(ram16sdp_inst_472_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(ram16sdp_inst_480_dout[2]),
  .I1(ram16sdp_inst_488_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(ram16sdp_inst_496_dout[2]),
  .I1(ram16sdp_inst_504_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(ram16sdp_inst_512_dout[2]),
  .I1(ram16sdp_inst_520_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(ram16sdp_inst_528_dout[2]),
  .I1(ram16sdp_inst_536_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(ram16sdp_inst_544_dout[2]),
  .I1(ram16sdp_inst_552_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(ram16sdp_inst_560_dout[2]),
  .I1(ram16sdp_inst_568_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(ram16sdp_inst_576_dout[2]),
  .I1(ram16sdp_inst_584_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(ram16sdp_inst_592_dout[2]),
  .I1(ram16sdp_inst_600_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(ram16sdp_inst_608_dout[2]),
  .I1(ram16sdp_inst_616_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(ram16sdp_inst_624_dout[2]),
  .I1(ram16sdp_inst_632_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(ram16sdp_inst_640_dout[2]),
  .I1(ram16sdp_inst_648_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(ram16sdp_inst_656_dout[2]),
  .I1(ram16sdp_inst_664_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(ram16sdp_inst_672_dout[2]),
  .I1(ram16sdp_inst_680_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(ram16sdp_inst_688_dout[2]),
  .I1(ram16sdp_inst_696_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(ram16sdp_inst_704_dout[2]),
  .I1(ram16sdp_inst_712_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(ram16sdp_inst_720_dout[2]),
  .I1(ram16sdp_inst_728_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(ram16sdp_inst_736_dout[2]),
  .I1(ram16sdp_inst_744_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(ram16sdp_inst_752_dout[2]),
  .I1(ram16sdp_inst_760_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(ram16sdp_inst_768_dout[2]),
  .I1(ram16sdp_inst_776_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(ram16sdp_inst_784_dout[2]),
  .I1(ram16sdp_inst_792_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(ram16sdp_inst_800_dout[2]),
  .I1(ram16sdp_inst_808_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(ram16sdp_inst_816_dout[2]),
  .I1(ram16sdp_inst_824_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(ram16sdp_inst_832_dout[2]),
  .I1(ram16sdp_inst_840_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(ram16sdp_inst_848_dout[2]),
  .I1(ram16sdp_inst_856_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(ram16sdp_inst_864_dout[2]),
  .I1(ram16sdp_inst_872_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(ram16sdp_inst_880_dout[2]),
  .I1(ram16sdp_inst_888_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(ram16sdp_inst_896_dout[2]),
  .I1(ram16sdp_inst_904_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(ram16sdp_inst_912_dout[2]),
  .I1(ram16sdp_inst_920_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(ram16sdp_inst_928_dout[2]),
  .I1(ram16sdp_inst_936_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(ram16sdp_inst_944_dout[2]),
  .I1(ram16sdp_inst_952_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_314 (
  .O(mux_o_314),
  .I0(ram16sdp_inst_960_dout[2]),
  .I1(ram16sdp_inst_968_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(ram16sdp_inst_976_dout[2]),
  .I1(ram16sdp_inst_984_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(ram16sdp_inst_992_dout[2]),
  .I1(ram16sdp_inst_1000_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(ram16sdp_inst_1008_dout[2]),
  .I1(ram16sdp_inst_1016_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(rad[5])
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(rad[5])
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(mux_o_258),
  .I1(mux_o_259),
  .S0(rad[5])
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(mux_o_260),
  .I1(mux_o_261),
  .S0(rad[5])
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(mux_o_262),
  .I1(mux_o_263),
  .S0(rad[5])
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(mux_o_264),
  .I1(mux_o_265),
  .S0(rad[5])
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(rad[5])
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(rad[5])
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(rad[5])
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(rad[5])
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(rad[5])
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(rad[5])
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(rad[5])
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(rad[5])
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(rad[5])
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(mux_o_284),
  .I1(mux_o_285),
  .S0(rad[5])
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(mux_o_286),
  .I1(mux_o_287),
  .S0(rad[5])
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(mux_o_288),
  .I1(mux_o_289),
  .S0(rad[5])
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(mux_o_290),
  .I1(mux_o_291),
  .S0(rad[5])
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(mux_o_292),
  .I1(mux_o_293),
  .S0(rad[5])
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_294),
  .I1(mux_o_295),
  .S0(rad[5])
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_296),
  .I1(mux_o_297),
  .S0(rad[5])
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(rad[5])
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(rad[5])
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(rad[5])
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(mux_o_304),
  .I1(mux_o_305),
  .S0(rad[5])
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(mux_o_306),
  .I1(mux_o_307),
  .S0(rad[5])
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(rad[5])
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(rad[5])
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(rad[5])
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_314),
  .I1(mux_o_315),
  .S0(rad[5])
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(mux_o_316),
  .I1(mux_o_317),
  .S0(rad[5])
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(mux_o_318),
  .I1(mux_o_319),
  .S0(rad[6])
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(mux_o_320),
  .I1(mux_o_321),
  .S0(rad[6])
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(rad[6])
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(rad[6])
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(rad[6])
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_328),
  .I1(mux_o_329),
  .S0(rad[6])
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(rad[6])
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(rad[6])
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(rad[6])
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(rad[6])
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(rad[6])
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(rad[6])
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_342),
  .I1(mux_o_343),
  .S0(rad[6])
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(mux_o_344),
  .I1(mux_o_345),
  .S0(rad[6])
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(mux_o_346),
  .I1(mux_o_347),
  .S0(rad[6])
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(mux_o_348),
  .I1(mux_o_349),
  .S0(rad[6])
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(rad[7])
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(rad[7])
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(rad[7])
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_356),
  .I1(mux_o_357),
  .S0(rad[7])
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_358),
  .I1(mux_o_359),
  .S0(rad[7])
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(mux_o_360),
  .I1(mux_o_361),
  .S0(rad[7])
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(mux_o_362),
  .I1(mux_o_363),
  .S0(rad[7])
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(rad[7])
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(rad[8])
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(rad[8])
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(mux_o_370),
  .I1(mux_o_371),
  .S0(rad[8])
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(rad[8])
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(mux_o_374),
  .I1(mux_o_375),
  .S0(rad[9])
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(mux_o_376),
  .I1(mux_o_377),
  .S0(rad[9])
);
MUX2 mux_inst_380 (
  .O(dout[2]),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(rad[10])
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(ram16sdp_inst_0_dout[3]),
  .I1(ram16sdp_inst_8_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(ram16sdp_inst_16_dout[3]),
  .I1(ram16sdp_inst_24_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(ram16sdp_inst_32_dout[3]),
  .I1(ram16sdp_inst_40_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(ram16sdp_inst_48_dout[3]),
  .I1(ram16sdp_inst_56_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(ram16sdp_inst_64_dout[3]),
  .I1(ram16sdp_inst_72_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(ram16sdp_inst_80_dout[3]),
  .I1(ram16sdp_inst_88_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(ram16sdp_inst_96_dout[3]),
  .I1(ram16sdp_inst_104_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(ram16sdp_inst_112_dout[3]),
  .I1(ram16sdp_inst_120_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(ram16sdp_inst_128_dout[3]),
  .I1(ram16sdp_inst_136_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(ram16sdp_inst_144_dout[3]),
  .I1(ram16sdp_inst_152_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(ram16sdp_inst_160_dout[3]),
  .I1(ram16sdp_inst_168_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(ram16sdp_inst_176_dout[3]),
  .I1(ram16sdp_inst_184_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(ram16sdp_inst_192_dout[3]),
  .I1(ram16sdp_inst_200_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(ram16sdp_inst_208_dout[3]),
  .I1(ram16sdp_inst_216_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(ram16sdp_inst_224_dout[3]),
  .I1(ram16sdp_inst_232_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(ram16sdp_inst_240_dout[3]),
  .I1(ram16sdp_inst_248_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(ram16sdp_inst_256_dout[3]),
  .I1(ram16sdp_inst_264_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(ram16sdp_inst_272_dout[3]),
  .I1(ram16sdp_inst_280_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(ram16sdp_inst_288_dout[3]),
  .I1(ram16sdp_inst_296_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(ram16sdp_inst_304_dout[3]),
  .I1(ram16sdp_inst_312_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(ram16sdp_inst_320_dout[3]),
  .I1(ram16sdp_inst_328_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(ram16sdp_inst_336_dout[3]),
  .I1(ram16sdp_inst_344_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(ram16sdp_inst_352_dout[3]),
  .I1(ram16sdp_inst_360_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(ram16sdp_inst_368_dout[3]),
  .I1(ram16sdp_inst_376_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(ram16sdp_inst_384_dout[3]),
  .I1(ram16sdp_inst_392_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(ram16sdp_inst_400_dout[3]),
  .I1(ram16sdp_inst_408_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(ram16sdp_inst_416_dout[3]),
  .I1(ram16sdp_inst_424_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(ram16sdp_inst_432_dout[3]),
  .I1(ram16sdp_inst_440_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(ram16sdp_inst_448_dout[3]),
  .I1(ram16sdp_inst_456_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(ram16sdp_inst_464_dout[3]),
  .I1(ram16sdp_inst_472_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(ram16sdp_inst_480_dout[3]),
  .I1(ram16sdp_inst_488_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(ram16sdp_inst_496_dout[3]),
  .I1(ram16sdp_inst_504_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(ram16sdp_inst_512_dout[3]),
  .I1(ram16sdp_inst_520_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(ram16sdp_inst_528_dout[3]),
  .I1(ram16sdp_inst_536_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(ram16sdp_inst_544_dout[3]),
  .I1(ram16sdp_inst_552_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(ram16sdp_inst_560_dout[3]),
  .I1(ram16sdp_inst_568_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(ram16sdp_inst_576_dout[3]),
  .I1(ram16sdp_inst_584_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(ram16sdp_inst_592_dout[3]),
  .I1(ram16sdp_inst_600_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_419 (
  .O(mux_o_419),
  .I0(ram16sdp_inst_608_dout[3]),
  .I1(ram16sdp_inst_616_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(ram16sdp_inst_624_dout[3]),
  .I1(ram16sdp_inst_632_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(ram16sdp_inst_640_dout[3]),
  .I1(ram16sdp_inst_648_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(ram16sdp_inst_656_dout[3]),
  .I1(ram16sdp_inst_664_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(ram16sdp_inst_672_dout[3]),
  .I1(ram16sdp_inst_680_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(ram16sdp_inst_688_dout[3]),
  .I1(ram16sdp_inst_696_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(ram16sdp_inst_704_dout[3]),
  .I1(ram16sdp_inst_712_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(ram16sdp_inst_720_dout[3]),
  .I1(ram16sdp_inst_728_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(ram16sdp_inst_736_dout[3]),
  .I1(ram16sdp_inst_744_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(ram16sdp_inst_752_dout[3]),
  .I1(ram16sdp_inst_760_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(ram16sdp_inst_768_dout[3]),
  .I1(ram16sdp_inst_776_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(ram16sdp_inst_784_dout[3]),
  .I1(ram16sdp_inst_792_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(ram16sdp_inst_800_dout[3]),
  .I1(ram16sdp_inst_808_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(ram16sdp_inst_816_dout[3]),
  .I1(ram16sdp_inst_824_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(ram16sdp_inst_832_dout[3]),
  .I1(ram16sdp_inst_840_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(ram16sdp_inst_848_dout[3]),
  .I1(ram16sdp_inst_856_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(ram16sdp_inst_864_dout[3]),
  .I1(ram16sdp_inst_872_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(ram16sdp_inst_880_dout[3]),
  .I1(ram16sdp_inst_888_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(ram16sdp_inst_896_dout[3]),
  .I1(ram16sdp_inst_904_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(ram16sdp_inst_912_dout[3]),
  .I1(ram16sdp_inst_920_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(ram16sdp_inst_928_dout[3]),
  .I1(ram16sdp_inst_936_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(ram16sdp_inst_944_dout[3]),
  .I1(ram16sdp_inst_952_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(ram16sdp_inst_960_dout[3]),
  .I1(ram16sdp_inst_968_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(ram16sdp_inst_976_dout[3]),
  .I1(ram16sdp_inst_984_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(ram16sdp_inst_992_dout[3]),
  .I1(ram16sdp_inst_1000_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(ram16sdp_inst_1008_dout[3]),
  .I1(ram16sdp_inst_1016_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(mux_o_381),
  .I1(mux_o_382),
  .S0(rad[5])
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(mux_o_383),
  .I1(mux_o_384),
  .S0(rad[5])
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(mux_o_385),
  .I1(mux_o_386),
  .S0(rad[5])
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(mux_o_387),
  .I1(mux_o_388),
  .S0(rad[5])
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(mux_o_389),
  .I1(mux_o_390),
  .S0(rad[5])
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(mux_o_391),
  .I1(mux_o_392),
  .S0(rad[5])
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(mux_o_393),
  .I1(mux_o_394),
  .S0(rad[5])
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(mux_o_395),
  .I1(mux_o_396),
  .S0(rad[5])
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(mux_o_397),
  .I1(mux_o_398),
  .S0(rad[5])
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(mux_o_399),
  .I1(mux_o_400),
  .S0(rad[5])
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(mux_o_401),
  .I1(mux_o_402),
  .S0(rad[5])
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_403),
  .I1(mux_o_404),
  .S0(rad[5])
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_405),
  .I1(mux_o_406),
  .S0(rad[5])
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_407),
  .I1(mux_o_408),
  .S0(rad[5])
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(rad[5])
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_411),
  .I1(mux_o_412),
  .S0(rad[5])
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(rad[5])
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_415),
  .I1(mux_o_416),
  .S0(rad[5])
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_417),
  .I1(mux_o_418),
  .S0(rad[5])
);
MUX2 mux_inst_464 (
  .O(mux_o_464),
  .I0(mux_o_419),
  .I1(mux_o_420),
  .S0(rad[5])
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(mux_o_421),
  .I1(mux_o_422),
  .S0(rad[5])
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(mux_o_423),
  .I1(mux_o_424),
  .S0(rad[5])
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(mux_o_425),
  .I1(mux_o_426),
  .S0(rad[5])
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(mux_o_427),
  .I1(mux_o_428),
  .S0(rad[5])
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(mux_o_429),
  .I1(mux_o_430),
  .S0(rad[5])
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(mux_o_431),
  .I1(mux_o_432),
  .S0(rad[5])
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(mux_o_433),
  .I1(mux_o_434),
  .S0(rad[5])
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(mux_o_435),
  .I1(mux_o_436),
  .S0(rad[5])
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_437),
  .I1(mux_o_438),
  .S0(rad[5])
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_439),
  .I1(mux_o_440),
  .S0(rad[5])
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(rad[5])
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(rad[5])
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(rad[6])
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(rad[6])
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(mux_o_449),
  .I1(mux_o_450),
  .S0(rad[6])
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(mux_o_451),
  .I1(mux_o_452),
  .S0(rad[6])
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(mux_o_453),
  .I1(mux_o_454),
  .S0(rad[6])
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(mux_o_455),
  .I1(mux_o_456),
  .S0(rad[6])
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(mux_o_457),
  .I1(mux_o_458),
  .S0(rad[6])
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(mux_o_459),
  .I1(mux_o_460),
  .S0(rad[6])
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(mux_o_461),
  .I1(mux_o_462),
  .S0(rad[6])
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(mux_o_463),
  .I1(mux_o_464),
  .S0(rad[6])
);
MUX2 mux_inst_487 (
  .O(mux_o_487),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(rad[6])
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(rad[6])
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(rad[6])
);
MUX2 mux_inst_490 (
  .O(mux_o_490),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(rad[6])
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(rad[6])
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(rad[6])
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(rad[7])
);
MUX2 mux_inst_494 (
  .O(mux_o_494),
  .I0(mux_o_479),
  .I1(mux_o_480),
  .S0(rad[7])
);
MUX2 mux_inst_495 (
  .O(mux_o_495),
  .I0(mux_o_481),
  .I1(mux_o_482),
  .S0(rad[7])
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(mux_o_483),
  .I1(mux_o_484),
  .S0(rad[7])
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(mux_o_485),
  .I1(mux_o_486),
  .S0(rad[7])
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(mux_o_487),
  .I1(mux_o_488),
  .S0(rad[7])
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(mux_o_489),
  .I1(mux_o_490),
  .S0(rad[7])
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(mux_o_491),
  .I1(mux_o_492),
  .S0(rad[7])
);
MUX2 mux_inst_501 (
  .O(mux_o_501),
  .I0(mux_o_493),
  .I1(mux_o_494),
  .S0(rad[8])
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(mux_o_495),
  .I1(mux_o_496),
  .S0(rad[8])
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(mux_o_497),
  .I1(mux_o_498),
  .S0(rad[8])
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(mux_o_499),
  .I1(mux_o_500),
  .S0(rad[8])
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(mux_o_501),
  .I1(mux_o_502),
  .S0(rad[9])
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(mux_o_503),
  .I1(mux_o_504),
  .S0(rad[9])
);
MUX2 mux_inst_507 (
  .O(dout[3]),
  .I0(mux_o_505),
  .I1(mux_o_506),
  .S0(rad[10])
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(ram16sdp_inst_1_dout[4]),
  .I1(ram16sdp_inst_9_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_509 (
  .O(mux_o_509),
  .I0(ram16sdp_inst_17_dout[4]),
  .I1(ram16sdp_inst_25_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(ram16sdp_inst_33_dout[4]),
  .I1(ram16sdp_inst_41_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(ram16sdp_inst_49_dout[4]),
  .I1(ram16sdp_inst_57_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(ram16sdp_inst_65_dout[4]),
  .I1(ram16sdp_inst_73_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(ram16sdp_inst_81_dout[4]),
  .I1(ram16sdp_inst_89_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(ram16sdp_inst_97_dout[4]),
  .I1(ram16sdp_inst_105_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_515 (
  .O(mux_o_515),
  .I0(ram16sdp_inst_113_dout[4]),
  .I1(ram16sdp_inst_121_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(ram16sdp_inst_129_dout[4]),
  .I1(ram16sdp_inst_137_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(ram16sdp_inst_145_dout[4]),
  .I1(ram16sdp_inst_153_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_518 (
  .O(mux_o_518),
  .I0(ram16sdp_inst_161_dout[4]),
  .I1(ram16sdp_inst_169_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(ram16sdp_inst_177_dout[4]),
  .I1(ram16sdp_inst_185_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(ram16sdp_inst_193_dout[4]),
  .I1(ram16sdp_inst_201_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(ram16sdp_inst_209_dout[4]),
  .I1(ram16sdp_inst_217_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(ram16sdp_inst_225_dout[4]),
  .I1(ram16sdp_inst_233_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(ram16sdp_inst_241_dout[4]),
  .I1(ram16sdp_inst_249_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_524 (
  .O(mux_o_524),
  .I0(ram16sdp_inst_257_dout[4]),
  .I1(ram16sdp_inst_265_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(ram16sdp_inst_273_dout[4]),
  .I1(ram16sdp_inst_281_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_526 (
  .O(mux_o_526),
  .I0(ram16sdp_inst_289_dout[4]),
  .I1(ram16sdp_inst_297_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(ram16sdp_inst_305_dout[4]),
  .I1(ram16sdp_inst_313_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(ram16sdp_inst_321_dout[4]),
  .I1(ram16sdp_inst_329_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_529 (
  .O(mux_o_529),
  .I0(ram16sdp_inst_337_dout[4]),
  .I1(ram16sdp_inst_345_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(ram16sdp_inst_353_dout[4]),
  .I1(ram16sdp_inst_361_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(ram16sdp_inst_369_dout[4]),
  .I1(ram16sdp_inst_377_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_532 (
  .O(mux_o_532),
  .I0(ram16sdp_inst_385_dout[4]),
  .I1(ram16sdp_inst_393_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(ram16sdp_inst_401_dout[4]),
  .I1(ram16sdp_inst_409_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(ram16sdp_inst_417_dout[4]),
  .I1(ram16sdp_inst_425_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(ram16sdp_inst_433_dout[4]),
  .I1(ram16sdp_inst_441_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(ram16sdp_inst_449_dout[4]),
  .I1(ram16sdp_inst_457_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(ram16sdp_inst_465_dout[4]),
  .I1(ram16sdp_inst_473_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(ram16sdp_inst_481_dout[4]),
  .I1(ram16sdp_inst_489_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_539 (
  .O(mux_o_539),
  .I0(ram16sdp_inst_497_dout[4]),
  .I1(ram16sdp_inst_505_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(ram16sdp_inst_513_dout[4]),
  .I1(ram16sdp_inst_521_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(ram16sdp_inst_529_dout[4]),
  .I1(ram16sdp_inst_537_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(ram16sdp_inst_545_dout[4]),
  .I1(ram16sdp_inst_553_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(ram16sdp_inst_561_dout[4]),
  .I1(ram16sdp_inst_569_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(ram16sdp_inst_577_dout[4]),
  .I1(ram16sdp_inst_585_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(ram16sdp_inst_593_dout[4]),
  .I1(ram16sdp_inst_601_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(ram16sdp_inst_609_dout[4]),
  .I1(ram16sdp_inst_617_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(ram16sdp_inst_625_dout[4]),
  .I1(ram16sdp_inst_633_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(ram16sdp_inst_641_dout[4]),
  .I1(ram16sdp_inst_649_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(ram16sdp_inst_657_dout[4]),
  .I1(ram16sdp_inst_665_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(ram16sdp_inst_673_dout[4]),
  .I1(ram16sdp_inst_681_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(ram16sdp_inst_689_dout[4]),
  .I1(ram16sdp_inst_697_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(ram16sdp_inst_705_dout[4]),
  .I1(ram16sdp_inst_713_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(ram16sdp_inst_721_dout[4]),
  .I1(ram16sdp_inst_729_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(ram16sdp_inst_737_dout[4]),
  .I1(ram16sdp_inst_745_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(ram16sdp_inst_753_dout[4]),
  .I1(ram16sdp_inst_761_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(ram16sdp_inst_769_dout[4]),
  .I1(ram16sdp_inst_777_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_557 (
  .O(mux_o_557),
  .I0(ram16sdp_inst_785_dout[4]),
  .I1(ram16sdp_inst_793_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(ram16sdp_inst_801_dout[4]),
  .I1(ram16sdp_inst_809_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(ram16sdp_inst_817_dout[4]),
  .I1(ram16sdp_inst_825_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(ram16sdp_inst_833_dout[4]),
  .I1(ram16sdp_inst_841_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(ram16sdp_inst_849_dout[4]),
  .I1(ram16sdp_inst_857_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(ram16sdp_inst_865_dout[4]),
  .I1(ram16sdp_inst_873_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(ram16sdp_inst_881_dout[4]),
  .I1(ram16sdp_inst_889_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(ram16sdp_inst_897_dout[4]),
  .I1(ram16sdp_inst_905_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(ram16sdp_inst_913_dout[4]),
  .I1(ram16sdp_inst_921_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_566 (
  .O(mux_o_566),
  .I0(ram16sdp_inst_929_dout[4]),
  .I1(ram16sdp_inst_937_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(ram16sdp_inst_945_dout[4]),
  .I1(ram16sdp_inst_953_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(ram16sdp_inst_961_dout[4]),
  .I1(ram16sdp_inst_969_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(ram16sdp_inst_977_dout[4]),
  .I1(ram16sdp_inst_985_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(ram16sdp_inst_993_dout[4]),
  .I1(ram16sdp_inst_1001_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_571 (
  .O(mux_o_571),
  .I0(ram16sdp_inst_1009_dout[4]),
  .I1(ram16sdp_inst_1017_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(mux_o_508),
  .I1(mux_o_509),
  .S0(rad[5])
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(mux_o_510),
  .I1(mux_o_511),
  .S0(rad[5])
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(rad[5])
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(mux_o_514),
  .I1(mux_o_515),
  .S0(rad[5])
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(rad[5])
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(mux_o_518),
  .I1(mux_o_519),
  .S0(rad[5])
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(mux_o_520),
  .I1(mux_o_521),
  .S0(rad[5])
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(rad[5])
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(mux_o_524),
  .I1(mux_o_525),
  .S0(rad[5])
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(mux_o_526),
  .I1(mux_o_527),
  .S0(rad[5])
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(mux_o_528),
  .I1(mux_o_529),
  .S0(rad[5])
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(mux_o_530),
  .I1(mux_o_531),
  .S0(rad[5])
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(mux_o_532),
  .I1(mux_o_533),
  .S0(rad[5])
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(mux_o_534),
  .I1(mux_o_535),
  .S0(rad[5])
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(mux_o_536),
  .I1(mux_o_537),
  .S0(rad[5])
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(mux_o_538),
  .I1(mux_o_539),
  .S0(rad[5])
);
MUX2 mux_inst_588 (
  .O(mux_o_588),
  .I0(mux_o_540),
  .I1(mux_o_541),
  .S0(rad[5])
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(mux_o_542),
  .I1(mux_o_543),
  .S0(rad[5])
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(mux_o_544),
  .I1(mux_o_545),
  .S0(rad[5])
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(mux_o_546),
  .I1(mux_o_547),
  .S0(rad[5])
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(mux_o_548),
  .I1(mux_o_549),
  .S0(rad[5])
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(mux_o_550),
  .I1(mux_o_551),
  .S0(rad[5])
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(mux_o_552),
  .I1(mux_o_553),
  .S0(rad[5])
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(mux_o_554),
  .I1(mux_o_555),
  .S0(rad[5])
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(mux_o_556),
  .I1(mux_o_557),
  .S0(rad[5])
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(mux_o_558),
  .I1(mux_o_559),
  .S0(rad[5])
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(rad[5])
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(mux_o_562),
  .I1(mux_o_563),
  .S0(rad[5])
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(mux_o_564),
  .I1(mux_o_565),
  .S0(rad[5])
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(mux_o_566),
  .I1(mux_o_567),
  .S0(rad[5])
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(mux_o_568),
  .I1(mux_o_569),
  .S0(rad[5])
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(mux_o_570),
  .I1(mux_o_571),
  .S0(rad[5])
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(mux_o_572),
  .I1(mux_o_573),
  .S0(rad[6])
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(mux_o_574),
  .I1(mux_o_575),
  .S0(rad[6])
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(mux_o_576),
  .I1(mux_o_577),
  .S0(rad[6])
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(mux_o_578),
  .I1(mux_o_579),
  .S0(rad[6])
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(mux_o_580),
  .I1(mux_o_581),
  .S0(rad[6])
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(mux_o_582),
  .I1(mux_o_583),
  .S0(rad[6])
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_584),
  .I1(mux_o_585),
  .S0(rad[6])
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_586),
  .I1(mux_o_587),
  .S0(rad[6])
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_588),
  .I1(mux_o_589),
  .S0(rad[6])
);
MUX2 mux_inst_613 (
  .O(mux_o_613),
  .I0(mux_o_590),
  .I1(mux_o_591),
  .S0(rad[6])
);
MUX2 mux_inst_614 (
  .O(mux_o_614),
  .I0(mux_o_592),
  .I1(mux_o_593),
  .S0(rad[6])
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(mux_o_594),
  .I1(mux_o_595),
  .S0(rad[6])
);
MUX2 mux_inst_616 (
  .O(mux_o_616),
  .I0(mux_o_596),
  .I1(mux_o_597),
  .S0(rad[6])
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(mux_o_598),
  .I1(mux_o_599),
  .S0(rad[6])
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(mux_o_600),
  .I1(mux_o_601),
  .S0(rad[6])
);
MUX2 mux_inst_619 (
  .O(mux_o_619),
  .I0(mux_o_602),
  .I1(mux_o_603),
  .S0(rad[6])
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(mux_o_604),
  .I1(mux_o_605),
  .S0(rad[7])
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(mux_o_606),
  .I1(mux_o_607),
  .S0(rad[7])
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(mux_o_608),
  .I1(mux_o_609),
  .S0(rad[7])
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(mux_o_610),
  .I1(mux_o_611),
  .S0(rad[7])
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(mux_o_612),
  .I1(mux_o_613),
  .S0(rad[7])
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(mux_o_614),
  .I1(mux_o_615),
  .S0(rad[7])
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(mux_o_616),
  .I1(mux_o_617),
  .S0(rad[7])
);
MUX2 mux_inst_627 (
  .O(mux_o_627),
  .I0(mux_o_618),
  .I1(mux_o_619),
  .S0(rad[7])
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(mux_o_620),
  .I1(mux_o_621),
  .S0(rad[8])
);
MUX2 mux_inst_629 (
  .O(mux_o_629),
  .I0(mux_o_622),
  .I1(mux_o_623),
  .S0(rad[8])
);
MUX2 mux_inst_630 (
  .O(mux_o_630),
  .I0(mux_o_624),
  .I1(mux_o_625),
  .S0(rad[8])
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(mux_o_626),
  .I1(mux_o_627),
  .S0(rad[8])
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(mux_o_628),
  .I1(mux_o_629),
  .S0(rad[9])
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(mux_o_630),
  .I1(mux_o_631),
  .S0(rad[9])
);
MUX2 mux_inst_634 (
  .O(dout[4]),
  .I0(mux_o_632),
  .I1(mux_o_633),
  .S0(rad[10])
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(ram16sdp_inst_1_dout[5]),
  .I1(ram16sdp_inst_9_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(ram16sdp_inst_17_dout[5]),
  .I1(ram16sdp_inst_25_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(ram16sdp_inst_33_dout[5]),
  .I1(ram16sdp_inst_41_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(ram16sdp_inst_49_dout[5]),
  .I1(ram16sdp_inst_57_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(ram16sdp_inst_65_dout[5]),
  .I1(ram16sdp_inst_73_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(ram16sdp_inst_81_dout[5]),
  .I1(ram16sdp_inst_89_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_641 (
  .O(mux_o_641),
  .I0(ram16sdp_inst_97_dout[5]),
  .I1(ram16sdp_inst_105_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(ram16sdp_inst_113_dout[5]),
  .I1(ram16sdp_inst_121_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(ram16sdp_inst_129_dout[5]),
  .I1(ram16sdp_inst_137_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_644 (
  .O(mux_o_644),
  .I0(ram16sdp_inst_145_dout[5]),
  .I1(ram16sdp_inst_153_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(ram16sdp_inst_161_dout[5]),
  .I1(ram16sdp_inst_169_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(ram16sdp_inst_177_dout[5]),
  .I1(ram16sdp_inst_185_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(ram16sdp_inst_193_dout[5]),
  .I1(ram16sdp_inst_201_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(ram16sdp_inst_209_dout[5]),
  .I1(ram16sdp_inst_217_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(ram16sdp_inst_225_dout[5]),
  .I1(ram16sdp_inst_233_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_650 (
  .O(mux_o_650),
  .I0(ram16sdp_inst_241_dout[5]),
  .I1(ram16sdp_inst_249_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(ram16sdp_inst_257_dout[5]),
  .I1(ram16sdp_inst_265_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(ram16sdp_inst_273_dout[5]),
  .I1(ram16sdp_inst_281_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(ram16sdp_inst_289_dout[5]),
  .I1(ram16sdp_inst_297_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(ram16sdp_inst_305_dout[5]),
  .I1(ram16sdp_inst_313_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_655 (
  .O(mux_o_655),
  .I0(ram16sdp_inst_321_dout[5]),
  .I1(ram16sdp_inst_329_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(ram16sdp_inst_337_dout[5]),
  .I1(ram16sdp_inst_345_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(ram16sdp_inst_353_dout[5]),
  .I1(ram16sdp_inst_361_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_658 (
  .O(mux_o_658),
  .I0(ram16sdp_inst_369_dout[5]),
  .I1(ram16sdp_inst_377_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_659 (
  .O(mux_o_659),
  .I0(ram16sdp_inst_385_dout[5]),
  .I1(ram16sdp_inst_393_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(ram16sdp_inst_401_dout[5]),
  .I1(ram16sdp_inst_409_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(ram16sdp_inst_417_dout[5]),
  .I1(ram16sdp_inst_425_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(ram16sdp_inst_433_dout[5]),
  .I1(ram16sdp_inst_441_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(ram16sdp_inst_449_dout[5]),
  .I1(ram16sdp_inst_457_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(ram16sdp_inst_465_dout[5]),
  .I1(ram16sdp_inst_473_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(ram16sdp_inst_481_dout[5]),
  .I1(ram16sdp_inst_489_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(ram16sdp_inst_497_dout[5]),
  .I1(ram16sdp_inst_505_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(ram16sdp_inst_513_dout[5]),
  .I1(ram16sdp_inst_521_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(ram16sdp_inst_529_dout[5]),
  .I1(ram16sdp_inst_537_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(ram16sdp_inst_545_dout[5]),
  .I1(ram16sdp_inst_553_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(ram16sdp_inst_561_dout[5]),
  .I1(ram16sdp_inst_569_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(ram16sdp_inst_577_dout[5]),
  .I1(ram16sdp_inst_585_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(ram16sdp_inst_593_dout[5]),
  .I1(ram16sdp_inst_601_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(ram16sdp_inst_609_dout[5]),
  .I1(ram16sdp_inst_617_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(ram16sdp_inst_625_dout[5]),
  .I1(ram16sdp_inst_633_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(ram16sdp_inst_641_dout[5]),
  .I1(ram16sdp_inst_649_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(ram16sdp_inst_657_dout[5]),
  .I1(ram16sdp_inst_665_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(ram16sdp_inst_673_dout[5]),
  .I1(ram16sdp_inst_681_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(ram16sdp_inst_689_dout[5]),
  .I1(ram16sdp_inst_697_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(ram16sdp_inst_705_dout[5]),
  .I1(ram16sdp_inst_713_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(ram16sdp_inst_721_dout[5]),
  .I1(ram16sdp_inst_729_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_681 (
  .O(mux_o_681),
  .I0(ram16sdp_inst_737_dout[5]),
  .I1(ram16sdp_inst_745_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(ram16sdp_inst_753_dout[5]),
  .I1(ram16sdp_inst_761_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(ram16sdp_inst_769_dout[5]),
  .I1(ram16sdp_inst_777_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(ram16sdp_inst_785_dout[5]),
  .I1(ram16sdp_inst_793_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(ram16sdp_inst_801_dout[5]),
  .I1(ram16sdp_inst_809_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(ram16sdp_inst_817_dout[5]),
  .I1(ram16sdp_inst_825_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(ram16sdp_inst_833_dout[5]),
  .I1(ram16sdp_inst_841_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(ram16sdp_inst_849_dout[5]),
  .I1(ram16sdp_inst_857_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(ram16sdp_inst_865_dout[5]),
  .I1(ram16sdp_inst_873_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(ram16sdp_inst_881_dout[5]),
  .I1(ram16sdp_inst_889_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(ram16sdp_inst_897_dout[5]),
  .I1(ram16sdp_inst_905_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_692 (
  .O(mux_o_692),
  .I0(ram16sdp_inst_913_dout[5]),
  .I1(ram16sdp_inst_921_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(ram16sdp_inst_929_dout[5]),
  .I1(ram16sdp_inst_937_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(ram16sdp_inst_945_dout[5]),
  .I1(ram16sdp_inst_953_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(ram16sdp_inst_961_dout[5]),
  .I1(ram16sdp_inst_969_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(ram16sdp_inst_977_dout[5]),
  .I1(ram16sdp_inst_985_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(ram16sdp_inst_993_dout[5]),
  .I1(ram16sdp_inst_1001_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(ram16sdp_inst_1009_dout[5]),
  .I1(ram16sdp_inst_1017_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(mux_o_635),
  .I1(mux_o_636),
  .S0(rad[5])
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(mux_o_637),
  .I1(mux_o_638),
  .S0(rad[5])
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(mux_o_639),
  .I1(mux_o_640),
  .S0(rad[5])
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(mux_o_641),
  .I1(mux_o_642),
  .S0(rad[5])
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(mux_o_643),
  .I1(mux_o_644),
  .S0(rad[5])
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(mux_o_645),
  .I1(mux_o_646),
  .S0(rad[5])
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(mux_o_647),
  .I1(mux_o_648),
  .S0(rad[5])
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(mux_o_649),
  .I1(mux_o_650),
  .S0(rad[5])
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(mux_o_651),
  .I1(mux_o_652),
  .S0(rad[5])
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(mux_o_653),
  .I1(mux_o_654),
  .S0(rad[5])
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(mux_o_655),
  .I1(mux_o_656),
  .S0(rad[5])
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(mux_o_657),
  .I1(mux_o_658),
  .S0(rad[5])
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(mux_o_659),
  .I1(mux_o_660),
  .S0(rad[5])
);
MUX2 mux_inst_712 (
  .O(mux_o_712),
  .I0(mux_o_661),
  .I1(mux_o_662),
  .S0(rad[5])
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(mux_o_663),
  .I1(mux_o_664),
  .S0(rad[5])
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(mux_o_665),
  .I1(mux_o_666),
  .S0(rad[5])
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(mux_o_667),
  .I1(mux_o_668),
  .S0(rad[5])
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(mux_o_669),
  .I1(mux_o_670),
  .S0(rad[5])
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(mux_o_671),
  .I1(mux_o_672),
  .S0(rad[5])
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(mux_o_673),
  .I1(mux_o_674),
  .S0(rad[5])
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(mux_o_675),
  .I1(mux_o_676),
  .S0(rad[5])
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(mux_o_677),
  .I1(mux_o_678),
  .S0(rad[5])
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(mux_o_679),
  .I1(mux_o_680),
  .S0(rad[5])
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(mux_o_681),
  .I1(mux_o_682),
  .S0(rad[5])
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(mux_o_683),
  .I1(mux_o_684),
  .S0(rad[5])
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(mux_o_685),
  .I1(mux_o_686),
  .S0(rad[5])
);
MUX2 mux_inst_725 (
  .O(mux_o_725),
  .I0(mux_o_687),
  .I1(mux_o_688),
  .S0(rad[5])
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(mux_o_689),
  .I1(mux_o_690),
  .S0(rad[5])
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(mux_o_691),
  .I1(mux_o_692),
  .S0(rad[5])
);
MUX2 mux_inst_728 (
  .O(mux_o_728),
  .I0(mux_o_693),
  .I1(mux_o_694),
  .S0(rad[5])
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(mux_o_695),
  .I1(mux_o_696),
  .S0(rad[5])
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(mux_o_697),
  .I1(mux_o_698),
  .S0(rad[5])
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(mux_o_699),
  .I1(mux_o_700),
  .S0(rad[6])
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(mux_o_701),
  .I1(mux_o_702),
  .S0(rad[6])
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(mux_o_703),
  .I1(mux_o_704),
  .S0(rad[6])
);
MUX2 mux_inst_734 (
  .O(mux_o_734),
  .I0(mux_o_705),
  .I1(mux_o_706),
  .S0(rad[6])
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(mux_o_707),
  .I1(mux_o_708),
  .S0(rad[6])
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(mux_o_709),
  .I1(mux_o_710),
  .S0(rad[6])
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(mux_o_711),
  .I1(mux_o_712),
  .S0(rad[6])
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(mux_o_713),
  .I1(mux_o_714),
  .S0(rad[6])
);
MUX2 mux_inst_739 (
  .O(mux_o_739),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(rad[6])
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(rad[6])
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(mux_o_719),
  .I1(mux_o_720),
  .S0(rad[6])
);
MUX2 mux_inst_742 (
  .O(mux_o_742),
  .I0(mux_o_721),
  .I1(mux_o_722),
  .S0(rad[6])
);
MUX2 mux_inst_743 (
  .O(mux_o_743),
  .I0(mux_o_723),
  .I1(mux_o_724),
  .S0(rad[6])
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(mux_o_725),
  .I1(mux_o_726),
  .S0(rad[6])
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(mux_o_727),
  .I1(mux_o_728),
  .S0(rad[6])
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(mux_o_729),
  .I1(mux_o_730),
  .S0(rad[6])
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(mux_o_731),
  .I1(mux_o_732),
  .S0(rad[7])
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(mux_o_733),
  .I1(mux_o_734),
  .S0(rad[7])
);
MUX2 mux_inst_749 (
  .O(mux_o_749),
  .I0(mux_o_735),
  .I1(mux_o_736),
  .S0(rad[7])
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(mux_o_737),
  .I1(mux_o_738),
  .S0(rad[7])
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(mux_o_739),
  .I1(mux_o_740),
  .S0(rad[7])
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(mux_o_741),
  .I1(mux_o_742),
  .S0(rad[7])
);
MUX2 mux_inst_753 (
  .O(mux_o_753),
  .I0(mux_o_743),
  .I1(mux_o_744),
  .S0(rad[7])
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(mux_o_745),
  .I1(mux_o_746),
  .S0(rad[7])
);
MUX2 mux_inst_755 (
  .O(mux_o_755),
  .I0(mux_o_747),
  .I1(mux_o_748),
  .S0(rad[8])
);
MUX2 mux_inst_756 (
  .O(mux_o_756),
  .I0(mux_o_749),
  .I1(mux_o_750),
  .S0(rad[8])
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(mux_o_751),
  .I1(mux_o_752),
  .S0(rad[8])
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(mux_o_753),
  .I1(mux_o_754),
  .S0(rad[8])
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(mux_o_755),
  .I1(mux_o_756),
  .S0(rad[9])
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(mux_o_757),
  .I1(mux_o_758),
  .S0(rad[9])
);
MUX2 mux_inst_761 (
  .O(dout[5]),
  .I0(mux_o_759),
  .I1(mux_o_760),
  .S0(rad[10])
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(ram16sdp_inst_1_dout[6]),
  .I1(ram16sdp_inst_9_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(ram16sdp_inst_17_dout[6]),
  .I1(ram16sdp_inst_25_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_764 (
  .O(mux_o_764),
  .I0(ram16sdp_inst_33_dout[6]),
  .I1(ram16sdp_inst_41_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(ram16sdp_inst_49_dout[6]),
  .I1(ram16sdp_inst_57_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(ram16sdp_inst_65_dout[6]),
  .I1(ram16sdp_inst_73_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_767 (
  .O(mux_o_767),
  .I0(ram16sdp_inst_81_dout[6]),
  .I1(ram16sdp_inst_89_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(ram16sdp_inst_97_dout[6]),
  .I1(ram16sdp_inst_105_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(ram16sdp_inst_113_dout[6]),
  .I1(ram16sdp_inst_121_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_770 (
  .O(mux_o_770),
  .I0(ram16sdp_inst_129_dout[6]),
  .I1(ram16sdp_inst_137_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(ram16sdp_inst_145_dout[6]),
  .I1(ram16sdp_inst_153_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(ram16sdp_inst_161_dout[6]),
  .I1(ram16sdp_inst_169_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(ram16sdp_inst_177_dout[6]),
  .I1(ram16sdp_inst_185_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_774 (
  .O(mux_o_774),
  .I0(ram16sdp_inst_193_dout[6]),
  .I1(ram16sdp_inst_201_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(ram16sdp_inst_209_dout[6]),
  .I1(ram16sdp_inst_217_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(ram16sdp_inst_225_dout[6]),
  .I1(ram16sdp_inst_233_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(ram16sdp_inst_241_dout[6]),
  .I1(ram16sdp_inst_249_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(ram16sdp_inst_257_dout[6]),
  .I1(ram16sdp_inst_265_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_779 (
  .O(mux_o_779),
  .I0(ram16sdp_inst_273_dout[6]),
  .I1(ram16sdp_inst_281_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(ram16sdp_inst_289_dout[6]),
  .I1(ram16sdp_inst_297_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_781 (
  .O(mux_o_781),
  .I0(ram16sdp_inst_305_dout[6]),
  .I1(ram16sdp_inst_313_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(ram16sdp_inst_321_dout[6]),
  .I1(ram16sdp_inst_329_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(ram16sdp_inst_337_dout[6]),
  .I1(ram16sdp_inst_345_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_784 (
  .O(mux_o_784),
  .I0(ram16sdp_inst_353_dout[6]),
  .I1(ram16sdp_inst_361_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(ram16sdp_inst_369_dout[6]),
  .I1(ram16sdp_inst_377_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(ram16sdp_inst_385_dout[6]),
  .I1(ram16sdp_inst_393_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(ram16sdp_inst_401_dout[6]),
  .I1(ram16sdp_inst_409_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(ram16sdp_inst_417_dout[6]),
  .I1(ram16sdp_inst_425_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(ram16sdp_inst_433_dout[6]),
  .I1(ram16sdp_inst_441_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(ram16sdp_inst_449_dout[6]),
  .I1(ram16sdp_inst_457_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(ram16sdp_inst_465_dout[6]),
  .I1(ram16sdp_inst_473_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(ram16sdp_inst_481_dout[6]),
  .I1(ram16sdp_inst_489_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(ram16sdp_inst_497_dout[6]),
  .I1(ram16sdp_inst_505_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_794 (
  .O(mux_o_794),
  .I0(ram16sdp_inst_513_dout[6]),
  .I1(ram16sdp_inst_521_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(ram16sdp_inst_529_dout[6]),
  .I1(ram16sdp_inst_537_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(ram16sdp_inst_545_dout[6]),
  .I1(ram16sdp_inst_553_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(ram16sdp_inst_561_dout[6]),
  .I1(ram16sdp_inst_569_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_798 (
  .O(mux_o_798),
  .I0(ram16sdp_inst_577_dout[6]),
  .I1(ram16sdp_inst_585_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(ram16sdp_inst_593_dout[6]),
  .I1(ram16sdp_inst_601_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(ram16sdp_inst_609_dout[6]),
  .I1(ram16sdp_inst_617_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_801 (
  .O(mux_o_801),
  .I0(ram16sdp_inst_625_dout[6]),
  .I1(ram16sdp_inst_633_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(ram16sdp_inst_641_dout[6]),
  .I1(ram16sdp_inst_649_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(ram16sdp_inst_657_dout[6]),
  .I1(ram16sdp_inst_665_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(ram16sdp_inst_673_dout[6]),
  .I1(ram16sdp_inst_681_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_805 (
  .O(mux_o_805),
  .I0(ram16sdp_inst_689_dout[6]),
  .I1(ram16sdp_inst_697_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(ram16sdp_inst_705_dout[6]),
  .I1(ram16sdp_inst_713_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(ram16sdp_inst_721_dout[6]),
  .I1(ram16sdp_inst_729_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(ram16sdp_inst_737_dout[6]),
  .I1(ram16sdp_inst_745_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_809 (
  .O(mux_o_809),
  .I0(ram16sdp_inst_753_dout[6]),
  .I1(ram16sdp_inst_761_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(ram16sdp_inst_769_dout[6]),
  .I1(ram16sdp_inst_777_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(ram16sdp_inst_785_dout[6]),
  .I1(ram16sdp_inst_793_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(ram16sdp_inst_801_dout[6]),
  .I1(ram16sdp_inst_809_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_813 (
  .O(mux_o_813),
  .I0(ram16sdp_inst_817_dout[6]),
  .I1(ram16sdp_inst_825_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_814 (
  .O(mux_o_814),
  .I0(ram16sdp_inst_833_dout[6]),
  .I1(ram16sdp_inst_841_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(ram16sdp_inst_849_dout[6]),
  .I1(ram16sdp_inst_857_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(ram16sdp_inst_865_dout[6]),
  .I1(ram16sdp_inst_873_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(ram16sdp_inst_881_dout[6]),
  .I1(ram16sdp_inst_889_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_818 (
  .O(mux_o_818),
  .I0(ram16sdp_inst_897_dout[6]),
  .I1(ram16sdp_inst_905_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(ram16sdp_inst_913_dout[6]),
  .I1(ram16sdp_inst_921_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(ram16sdp_inst_929_dout[6]),
  .I1(ram16sdp_inst_937_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(ram16sdp_inst_945_dout[6]),
  .I1(ram16sdp_inst_953_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(ram16sdp_inst_961_dout[6]),
  .I1(ram16sdp_inst_969_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(ram16sdp_inst_977_dout[6]),
  .I1(ram16sdp_inst_985_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(ram16sdp_inst_993_dout[6]),
  .I1(ram16sdp_inst_1001_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(ram16sdp_inst_1009_dout[6]),
  .I1(ram16sdp_inst_1017_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(mux_o_762),
  .I1(mux_o_763),
  .S0(rad[5])
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(mux_o_764),
  .I1(mux_o_765),
  .S0(rad[5])
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(mux_o_766),
  .I1(mux_o_767),
  .S0(rad[5])
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(mux_o_768),
  .I1(mux_o_769),
  .S0(rad[5])
);
MUX2 mux_inst_830 (
  .O(mux_o_830),
  .I0(mux_o_770),
  .I1(mux_o_771),
  .S0(rad[5])
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(mux_o_772),
  .I1(mux_o_773),
  .S0(rad[5])
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(mux_o_774),
  .I1(mux_o_775),
  .S0(rad[5])
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(mux_o_776),
  .I1(mux_o_777),
  .S0(rad[5])
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(mux_o_778),
  .I1(mux_o_779),
  .S0(rad[5])
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(mux_o_780),
  .I1(mux_o_781),
  .S0(rad[5])
);
MUX2 mux_inst_836 (
  .O(mux_o_836),
  .I0(mux_o_782),
  .I1(mux_o_783),
  .S0(rad[5])
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(mux_o_784),
  .I1(mux_o_785),
  .S0(rad[5])
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(mux_o_786),
  .I1(mux_o_787),
  .S0(rad[5])
);
MUX2 mux_inst_839 (
  .O(mux_o_839),
  .I0(mux_o_788),
  .I1(mux_o_789),
  .S0(rad[5])
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(mux_o_790),
  .I1(mux_o_791),
  .S0(rad[5])
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(mux_o_792),
  .I1(mux_o_793),
  .S0(rad[5])
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(mux_o_794),
  .I1(mux_o_795),
  .S0(rad[5])
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(mux_o_796),
  .I1(mux_o_797),
  .S0(rad[5])
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(mux_o_798),
  .I1(mux_o_799),
  .S0(rad[5])
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(mux_o_800),
  .I1(mux_o_801),
  .S0(rad[5])
);
MUX2 mux_inst_846 (
  .O(mux_o_846),
  .I0(mux_o_802),
  .I1(mux_o_803),
  .S0(rad[5])
);
MUX2 mux_inst_847 (
  .O(mux_o_847),
  .I0(mux_o_804),
  .I1(mux_o_805),
  .S0(rad[5])
);
MUX2 mux_inst_848 (
  .O(mux_o_848),
  .I0(mux_o_806),
  .I1(mux_o_807),
  .S0(rad[5])
);
MUX2 mux_inst_849 (
  .O(mux_o_849),
  .I0(mux_o_808),
  .I1(mux_o_809),
  .S0(rad[5])
);
MUX2 mux_inst_850 (
  .O(mux_o_850),
  .I0(mux_o_810),
  .I1(mux_o_811),
  .S0(rad[5])
);
MUX2 mux_inst_851 (
  .O(mux_o_851),
  .I0(mux_o_812),
  .I1(mux_o_813),
  .S0(rad[5])
);
MUX2 mux_inst_852 (
  .O(mux_o_852),
  .I0(mux_o_814),
  .I1(mux_o_815),
  .S0(rad[5])
);
MUX2 mux_inst_853 (
  .O(mux_o_853),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(rad[5])
);
MUX2 mux_inst_854 (
  .O(mux_o_854),
  .I0(mux_o_818),
  .I1(mux_o_819),
  .S0(rad[5])
);
MUX2 mux_inst_855 (
  .O(mux_o_855),
  .I0(mux_o_820),
  .I1(mux_o_821),
  .S0(rad[5])
);
MUX2 mux_inst_856 (
  .O(mux_o_856),
  .I0(mux_o_822),
  .I1(mux_o_823),
  .S0(rad[5])
);
MUX2 mux_inst_857 (
  .O(mux_o_857),
  .I0(mux_o_824),
  .I1(mux_o_825),
  .S0(rad[5])
);
MUX2 mux_inst_858 (
  .O(mux_o_858),
  .I0(mux_o_826),
  .I1(mux_o_827),
  .S0(rad[6])
);
MUX2 mux_inst_859 (
  .O(mux_o_859),
  .I0(mux_o_828),
  .I1(mux_o_829),
  .S0(rad[6])
);
MUX2 mux_inst_860 (
  .O(mux_o_860),
  .I0(mux_o_830),
  .I1(mux_o_831),
  .S0(rad[6])
);
MUX2 mux_inst_861 (
  .O(mux_o_861),
  .I0(mux_o_832),
  .I1(mux_o_833),
  .S0(rad[6])
);
MUX2 mux_inst_862 (
  .O(mux_o_862),
  .I0(mux_o_834),
  .I1(mux_o_835),
  .S0(rad[6])
);
MUX2 mux_inst_863 (
  .O(mux_o_863),
  .I0(mux_o_836),
  .I1(mux_o_837),
  .S0(rad[6])
);
MUX2 mux_inst_864 (
  .O(mux_o_864),
  .I0(mux_o_838),
  .I1(mux_o_839),
  .S0(rad[6])
);
MUX2 mux_inst_865 (
  .O(mux_o_865),
  .I0(mux_o_840),
  .I1(mux_o_841),
  .S0(rad[6])
);
MUX2 mux_inst_866 (
  .O(mux_o_866),
  .I0(mux_o_842),
  .I1(mux_o_843),
  .S0(rad[6])
);
MUX2 mux_inst_867 (
  .O(mux_o_867),
  .I0(mux_o_844),
  .I1(mux_o_845),
  .S0(rad[6])
);
MUX2 mux_inst_868 (
  .O(mux_o_868),
  .I0(mux_o_846),
  .I1(mux_o_847),
  .S0(rad[6])
);
MUX2 mux_inst_869 (
  .O(mux_o_869),
  .I0(mux_o_848),
  .I1(mux_o_849),
  .S0(rad[6])
);
MUX2 mux_inst_870 (
  .O(mux_o_870),
  .I0(mux_o_850),
  .I1(mux_o_851),
  .S0(rad[6])
);
MUX2 mux_inst_871 (
  .O(mux_o_871),
  .I0(mux_o_852),
  .I1(mux_o_853),
  .S0(rad[6])
);
MUX2 mux_inst_872 (
  .O(mux_o_872),
  .I0(mux_o_854),
  .I1(mux_o_855),
  .S0(rad[6])
);
MUX2 mux_inst_873 (
  .O(mux_o_873),
  .I0(mux_o_856),
  .I1(mux_o_857),
  .S0(rad[6])
);
MUX2 mux_inst_874 (
  .O(mux_o_874),
  .I0(mux_o_858),
  .I1(mux_o_859),
  .S0(rad[7])
);
MUX2 mux_inst_875 (
  .O(mux_o_875),
  .I0(mux_o_860),
  .I1(mux_o_861),
  .S0(rad[7])
);
MUX2 mux_inst_876 (
  .O(mux_o_876),
  .I0(mux_o_862),
  .I1(mux_o_863),
  .S0(rad[7])
);
MUX2 mux_inst_877 (
  .O(mux_o_877),
  .I0(mux_o_864),
  .I1(mux_o_865),
  .S0(rad[7])
);
MUX2 mux_inst_878 (
  .O(mux_o_878),
  .I0(mux_o_866),
  .I1(mux_o_867),
  .S0(rad[7])
);
MUX2 mux_inst_879 (
  .O(mux_o_879),
  .I0(mux_o_868),
  .I1(mux_o_869),
  .S0(rad[7])
);
MUX2 mux_inst_880 (
  .O(mux_o_880),
  .I0(mux_o_870),
  .I1(mux_o_871),
  .S0(rad[7])
);
MUX2 mux_inst_881 (
  .O(mux_o_881),
  .I0(mux_o_872),
  .I1(mux_o_873),
  .S0(rad[7])
);
MUX2 mux_inst_882 (
  .O(mux_o_882),
  .I0(mux_o_874),
  .I1(mux_o_875),
  .S0(rad[8])
);
MUX2 mux_inst_883 (
  .O(mux_o_883),
  .I0(mux_o_876),
  .I1(mux_o_877),
  .S0(rad[8])
);
MUX2 mux_inst_884 (
  .O(mux_o_884),
  .I0(mux_o_878),
  .I1(mux_o_879),
  .S0(rad[8])
);
MUX2 mux_inst_885 (
  .O(mux_o_885),
  .I0(mux_o_880),
  .I1(mux_o_881),
  .S0(rad[8])
);
MUX2 mux_inst_886 (
  .O(mux_o_886),
  .I0(mux_o_882),
  .I1(mux_o_883),
  .S0(rad[9])
);
MUX2 mux_inst_887 (
  .O(mux_o_887),
  .I0(mux_o_884),
  .I1(mux_o_885),
  .S0(rad[9])
);
MUX2 mux_inst_888 (
  .O(dout[6]),
  .I0(mux_o_886),
  .I1(mux_o_887),
  .S0(rad[10])
);
MUX2 mux_inst_889 (
  .O(mux_o_889),
  .I0(ram16sdp_inst_1_dout[7]),
  .I1(ram16sdp_inst_9_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_890 (
  .O(mux_o_890),
  .I0(ram16sdp_inst_17_dout[7]),
  .I1(ram16sdp_inst_25_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_891 (
  .O(mux_o_891),
  .I0(ram16sdp_inst_33_dout[7]),
  .I1(ram16sdp_inst_41_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_892 (
  .O(mux_o_892),
  .I0(ram16sdp_inst_49_dout[7]),
  .I1(ram16sdp_inst_57_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_893 (
  .O(mux_o_893),
  .I0(ram16sdp_inst_65_dout[7]),
  .I1(ram16sdp_inst_73_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_894 (
  .O(mux_o_894),
  .I0(ram16sdp_inst_81_dout[7]),
  .I1(ram16sdp_inst_89_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_895 (
  .O(mux_o_895),
  .I0(ram16sdp_inst_97_dout[7]),
  .I1(ram16sdp_inst_105_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_896 (
  .O(mux_o_896),
  .I0(ram16sdp_inst_113_dout[7]),
  .I1(ram16sdp_inst_121_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_897 (
  .O(mux_o_897),
  .I0(ram16sdp_inst_129_dout[7]),
  .I1(ram16sdp_inst_137_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_898 (
  .O(mux_o_898),
  .I0(ram16sdp_inst_145_dout[7]),
  .I1(ram16sdp_inst_153_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_899 (
  .O(mux_o_899),
  .I0(ram16sdp_inst_161_dout[7]),
  .I1(ram16sdp_inst_169_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_900 (
  .O(mux_o_900),
  .I0(ram16sdp_inst_177_dout[7]),
  .I1(ram16sdp_inst_185_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_901 (
  .O(mux_o_901),
  .I0(ram16sdp_inst_193_dout[7]),
  .I1(ram16sdp_inst_201_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_902 (
  .O(mux_o_902),
  .I0(ram16sdp_inst_209_dout[7]),
  .I1(ram16sdp_inst_217_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_903 (
  .O(mux_o_903),
  .I0(ram16sdp_inst_225_dout[7]),
  .I1(ram16sdp_inst_233_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_904 (
  .O(mux_o_904),
  .I0(ram16sdp_inst_241_dout[7]),
  .I1(ram16sdp_inst_249_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_905 (
  .O(mux_o_905),
  .I0(ram16sdp_inst_257_dout[7]),
  .I1(ram16sdp_inst_265_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(ram16sdp_inst_273_dout[7]),
  .I1(ram16sdp_inst_281_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(ram16sdp_inst_289_dout[7]),
  .I1(ram16sdp_inst_297_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(ram16sdp_inst_305_dout[7]),
  .I1(ram16sdp_inst_313_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(ram16sdp_inst_321_dout[7]),
  .I1(ram16sdp_inst_329_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(ram16sdp_inst_337_dout[7]),
  .I1(ram16sdp_inst_345_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(ram16sdp_inst_353_dout[7]),
  .I1(ram16sdp_inst_361_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(ram16sdp_inst_369_dout[7]),
  .I1(ram16sdp_inst_377_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(ram16sdp_inst_385_dout[7]),
  .I1(ram16sdp_inst_393_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_914 (
  .O(mux_o_914),
  .I0(ram16sdp_inst_401_dout[7]),
  .I1(ram16sdp_inst_409_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(ram16sdp_inst_417_dout[7]),
  .I1(ram16sdp_inst_425_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(ram16sdp_inst_433_dout[7]),
  .I1(ram16sdp_inst_441_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(ram16sdp_inst_449_dout[7]),
  .I1(ram16sdp_inst_457_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(ram16sdp_inst_465_dout[7]),
  .I1(ram16sdp_inst_473_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(ram16sdp_inst_481_dout[7]),
  .I1(ram16sdp_inst_489_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(ram16sdp_inst_497_dout[7]),
  .I1(ram16sdp_inst_505_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(ram16sdp_inst_513_dout[7]),
  .I1(ram16sdp_inst_521_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(ram16sdp_inst_529_dout[7]),
  .I1(ram16sdp_inst_537_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(ram16sdp_inst_545_dout[7]),
  .I1(ram16sdp_inst_553_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(ram16sdp_inst_561_dout[7]),
  .I1(ram16sdp_inst_569_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(ram16sdp_inst_577_dout[7]),
  .I1(ram16sdp_inst_585_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(ram16sdp_inst_593_dout[7]),
  .I1(ram16sdp_inst_601_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(ram16sdp_inst_609_dout[7]),
  .I1(ram16sdp_inst_617_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(ram16sdp_inst_625_dout[7]),
  .I1(ram16sdp_inst_633_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_929 (
  .O(mux_o_929),
  .I0(ram16sdp_inst_641_dout[7]),
  .I1(ram16sdp_inst_649_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(ram16sdp_inst_657_dout[7]),
  .I1(ram16sdp_inst_665_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(ram16sdp_inst_673_dout[7]),
  .I1(ram16sdp_inst_681_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(ram16sdp_inst_689_dout[7]),
  .I1(ram16sdp_inst_697_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(ram16sdp_inst_705_dout[7]),
  .I1(ram16sdp_inst_713_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_934 (
  .O(mux_o_934),
  .I0(ram16sdp_inst_721_dout[7]),
  .I1(ram16sdp_inst_729_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_935 (
  .O(mux_o_935),
  .I0(ram16sdp_inst_737_dout[7]),
  .I1(ram16sdp_inst_745_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_936 (
  .O(mux_o_936),
  .I0(ram16sdp_inst_753_dout[7]),
  .I1(ram16sdp_inst_761_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(ram16sdp_inst_769_dout[7]),
  .I1(ram16sdp_inst_777_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(ram16sdp_inst_785_dout[7]),
  .I1(ram16sdp_inst_793_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(ram16sdp_inst_801_dout[7]),
  .I1(ram16sdp_inst_809_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(ram16sdp_inst_817_dout[7]),
  .I1(ram16sdp_inst_825_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(ram16sdp_inst_833_dout[7]),
  .I1(ram16sdp_inst_841_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(ram16sdp_inst_849_dout[7]),
  .I1(ram16sdp_inst_857_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(ram16sdp_inst_865_dout[7]),
  .I1(ram16sdp_inst_873_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_944 (
  .O(mux_o_944),
  .I0(ram16sdp_inst_881_dout[7]),
  .I1(ram16sdp_inst_889_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(ram16sdp_inst_897_dout[7]),
  .I1(ram16sdp_inst_905_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(ram16sdp_inst_913_dout[7]),
  .I1(ram16sdp_inst_921_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(ram16sdp_inst_929_dout[7]),
  .I1(ram16sdp_inst_937_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(ram16sdp_inst_945_dout[7]),
  .I1(ram16sdp_inst_953_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(ram16sdp_inst_961_dout[7]),
  .I1(ram16sdp_inst_969_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(ram16sdp_inst_977_dout[7]),
  .I1(ram16sdp_inst_985_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_951 (
  .O(mux_o_951),
  .I0(ram16sdp_inst_993_dout[7]),
  .I1(ram16sdp_inst_1001_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(ram16sdp_inst_1009_dout[7]),
  .I1(ram16sdp_inst_1017_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(mux_o_889),
  .I1(mux_o_890),
  .S0(rad[5])
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(mux_o_891),
  .I1(mux_o_892),
  .S0(rad[5])
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(mux_o_893),
  .I1(mux_o_894),
  .S0(rad[5])
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(mux_o_895),
  .I1(mux_o_896),
  .S0(rad[5])
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(mux_o_897),
  .I1(mux_o_898),
  .S0(rad[5])
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(mux_o_899),
  .I1(mux_o_900),
  .S0(rad[5])
);
MUX2 mux_inst_959 (
  .O(mux_o_959),
  .I0(mux_o_901),
  .I1(mux_o_902),
  .S0(rad[5])
);
MUX2 mux_inst_960 (
  .O(mux_o_960),
  .I0(mux_o_903),
  .I1(mux_o_904),
  .S0(rad[5])
);
MUX2 mux_inst_961 (
  .O(mux_o_961),
  .I0(mux_o_905),
  .I1(mux_o_906),
  .S0(rad[5])
);
MUX2 mux_inst_962 (
  .O(mux_o_962),
  .I0(mux_o_907),
  .I1(mux_o_908),
  .S0(rad[5])
);
MUX2 mux_inst_963 (
  .O(mux_o_963),
  .I0(mux_o_909),
  .I1(mux_o_910),
  .S0(rad[5])
);
MUX2 mux_inst_964 (
  .O(mux_o_964),
  .I0(mux_o_911),
  .I1(mux_o_912),
  .S0(rad[5])
);
MUX2 mux_inst_965 (
  .O(mux_o_965),
  .I0(mux_o_913),
  .I1(mux_o_914),
  .S0(rad[5])
);
MUX2 mux_inst_966 (
  .O(mux_o_966),
  .I0(mux_o_915),
  .I1(mux_o_916),
  .S0(rad[5])
);
MUX2 mux_inst_967 (
  .O(mux_o_967),
  .I0(mux_o_917),
  .I1(mux_o_918),
  .S0(rad[5])
);
MUX2 mux_inst_968 (
  .O(mux_o_968),
  .I0(mux_o_919),
  .I1(mux_o_920),
  .S0(rad[5])
);
MUX2 mux_inst_969 (
  .O(mux_o_969),
  .I0(mux_o_921),
  .I1(mux_o_922),
  .S0(rad[5])
);
MUX2 mux_inst_970 (
  .O(mux_o_970),
  .I0(mux_o_923),
  .I1(mux_o_924),
  .S0(rad[5])
);
MUX2 mux_inst_971 (
  .O(mux_o_971),
  .I0(mux_o_925),
  .I1(mux_o_926),
  .S0(rad[5])
);
MUX2 mux_inst_972 (
  .O(mux_o_972),
  .I0(mux_o_927),
  .I1(mux_o_928),
  .S0(rad[5])
);
MUX2 mux_inst_973 (
  .O(mux_o_973),
  .I0(mux_o_929),
  .I1(mux_o_930),
  .S0(rad[5])
);
MUX2 mux_inst_974 (
  .O(mux_o_974),
  .I0(mux_o_931),
  .I1(mux_o_932),
  .S0(rad[5])
);
MUX2 mux_inst_975 (
  .O(mux_o_975),
  .I0(mux_o_933),
  .I1(mux_o_934),
  .S0(rad[5])
);
MUX2 mux_inst_976 (
  .O(mux_o_976),
  .I0(mux_o_935),
  .I1(mux_o_936),
  .S0(rad[5])
);
MUX2 mux_inst_977 (
  .O(mux_o_977),
  .I0(mux_o_937),
  .I1(mux_o_938),
  .S0(rad[5])
);
MUX2 mux_inst_978 (
  .O(mux_o_978),
  .I0(mux_o_939),
  .I1(mux_o_940),
  .S0(rad[5])
);
MUX2 mux_inst_979 (
  .O(mux_o_979),
  .I0(mux_o_941),
  .I1(mux_o_942),
  .S0(rad[5])
);
MUX2 mux_inst_980 (
  .O(mux_o_980),
  .I0(mux_o_943),
  .I1(mux_o_944),
  .S0(rad[5])
);
MUX2 mux_inst_981 (
  .O(mux_o_981),
  .I0(mux_o_945),
  .I1(mux_o_946),
  .S0(rad[5])
);
MUX2 mux_inst_982 (
  .O(mux_o_982),
  .I0(mux_o_947),
  .I1(mux_o_948),
  .S0(rad[5])
);
MUX2 mux_inst_983 (
  .O(mux_o_983),
  .I0(mux_o_949),
  .I1(mux_o_950),
  .S0(rad[5])
);
MUX2 mux_inst_984 (
  .O(mux_o_984),
  .I0(mux_o_951),
  .I1(mux_o_952),
  .S0(rad[5])
);
MUX2 mux_inst_985 (
  .O(mux_o_985),
  .I0(mux_o_953),
  .I1(mux_o_954),
  .S0(rad[6])
);
MUX2 mux_inst_986 (
  .O(mux_o_986),
  .I0(mux_o_955),
  .I1(mux_o_956),
  .S0(rad[6])
);
MUX2 mux_inst_987 (
  .O(mux_o_987),
  .I0(mux_o_957),
  .I1(mux_o_958),
  .S0(rad[6])
);
MUX2 mux_inst_988 (
  .O(mux_o_988),
  .I0(mux_o_959),
  .I1(mux_o_960),
  .S0(rad[6])
);
MUX2 mux_inst_989 (
  .O(mux_o_989),
  .I0(mux_o_961),
  .I1(mux_o_962),
  .S0(rad[6])
);
MUX2 mux_inst_990 (
  .O(mux_o_990),
  .I0(mux_o_963),
  .I1(mux_o_964),
  .S0(rad[6])
);
MUX2 mux_inst_991 (
  .O(mux_o_991),
  .I0(mux_o_965),
  .I1(mux_o_966),
  .S0(rad[6])
);
MUX2 mux_inst_992 (
  .O(mux_o_992),
  .I0(mux_o_967),
  .I1(mux_o_968),
  .S0(rad[6])
);
MUX2 mux_inst_993 (
  .O(mux_o_993),
  .I0(mux_o_969),
  .I1(mux_o_970),
  .S0(rad[6])
);
MUX2 mux_inst_994 (
  .O(mux_o_994),
  .I0(mux_o_971),
  .I1(mux_o_972),
  .S0(rad[6])
);
MUX2 mux_inst_995 (
  .O(mux_o_995),
  .I0(mux_o_973),
  .I1(mux_o_974),
  .S0(rad[6])
);
MUX2 mux_inst_996 (
  .O(mux_o_996),
  .I0(mux_o_975),
  .I1(mux_o_976),
  .S0(rad[6])
);
MUX2 mux_inst_997 (
  .O(mux_o_997),
  .I0(mux_o_977),
  .I1(mux_o_978),
  .S0(rad[6])
);
MUX2 mux_inst_998 (
  .O(mux_o_998),
  .I0(mux_o_979),
  .I1(mux_o_980),
  .S0(rad[6])
);
MUX2 mux_inst_999 (
  .O(mux_o_999),
  .I0(mux_o_981),
  .I1(mux_o_982),
  .S0(rad[6])
);
MUX2 mux_inst_1000 (
  .O(mux_o_1000),
  .I0(mux_o_983),
  .I1(mux_o_984),
  .S0(rad[6])
);
MUX2 mux_inst_1001 (
  .O(mux_o_1001),
  .I0(mux_o_985),
  .I1(mux_o_986),
  .S0(rad[7])
);
MUX2 mux_inst_1002 (
  .O(mux_o_1002),
  .I0(mux_o_987),
  .I1(mux_o_988),
  .S0(rad[7])
);
MUX2 mux_inst_1003 (
  .O(mux_o_1003),
  .I0(mux_o_989),
  .I1(mux_o_990),
  .S0(rad[7])
);
MUX2 mux_inst_1004 (
  .O(mux_o_1004),
  .I0(mux_o_991),
  .I1(mux_o_992),
  .S0(rad[7])
);
MUX2 mux_inst_1005 (
  .O(mux_o_1005),
  .I0(mux_o_993),
  .I1(mux_o_994),
  .S0(rad[7])
);
MUX2 mux_inst_1006 (
  .O(mux_o_1006),
  .I0(mux_o_995),
  .I1(mux_o_996),
  .S0(rad[7])
);
MUX2 mux_inst_1007 (
  .O(mux_o_1007),
  .I0(mux_o_997),
  .I1(mux_o_998),
  .S0(rad[7])
);
MUX2 mux_inst_1008 (
  .O(mux_o_1008),
  .I0(mux_o_999),
  .I1(mux_o_1000),
  .S0(rad[7])
);
MUX2 mux_inst_1009 (
  .O(mux_o_1009),
  .I0(mux_o_1001),
  .I1(mux_o_1002),
  .S0(rad[8])
);
MUX2 mux_inst_1010 (
  .O(mux_o_1010),
  .I0(mux_o_1003),
  .I1(mux_o_1004),
  .S0(rad[8])
);
MUX2 mux_inst_1011 (
  .O(mux_o_1011),
  .I0(mux_o_1005),
  .I1(mux_o_1006),
  .S0(rad[8])
);
MUX2 mux_inst_1012 (
  .O(mux_o_1012),
  .I0(mux_o_1007),
  .I1(mux_o_1008),
  .S0(rad[8])
);
MUX2 mux_inst_1013 (
  .O(mux_o_1013),
  .I0(mux_o_1009),
  .I1(mux_o_1010),
  .S0(rad[9])
);
MUX2 mux_inst_1014 (
  .O(mux_o_1014),
  .I0(mux_o_1011),
  .I1(mux_o_1012),
  .S0(rad[9])
);
MUX2 mux_inst_1015 (
  .O(dout[7]),
  .I0(mux_o_1013),
  .I1(mux_o_1014),
  .S0(rad[10])
);
MUX2 mux_inst_1016 (
  .O(mux_o_1016),
  .I0(ram16sdp_inst_2_dout[8]),
  .I1(ram16sdp_inst_10_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1017 (
  .O(mux_o_1017),
  .I0(ram16sdp_inst_18_dout[8]),
  .I1(ram16sdp_inst_26_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1018 (
  .O(mux_o_1018),
  .I0(ram16sdp_inst_34_dout[8]),
  .I1(ram16sdp_inst_42_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1019 (
  .O(mux_o_1019),
  .I0(ram16sdp_inst_50_dout[8]),
  .I1(ram16sdp_inst_58_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1020 (
  .O(mux_o_1020),
  .I0(ram16sdp_inst_66_dout[8]),
  .I1(ram16sdp_inst_74_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1021 (
  .O(mux_o_1021),
  .I0(ram16sdp_inst_82_dout[8]),
  .I1(ram16sdp_inst_90_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1022 (
  .O(mux_o_1022),
  .I0(ram16sdp_inst_98_dout[8]),
  .I1(ram16sdp_inst_106_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1023 (
  .O(mux_o_1023),
  .I0(ram16sdp_inst_114_dout[8]),
  .I1(ram16sdp_inst_122_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1024 (
  .O(mux_o_1024),
  .I0(ram16sdp_inst_130_dout[8]),
  .I1(ram16sdp_inst_138_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1025 (
  .O(mux_o_1025),
  .I0(ram16sdp_inst_146_dout[8]),
  .I1(ram16sdp_inst_154_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1026 (
  .O(mux_o_1026),
  .I0(ram16sdp_inst_162_dout[8]),
  .I1(ram16sdp_inst_170_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1027 (
  .O(mux_o_1027),
  .I0(ram16sdp_inst_178_dout[8]),
  .I1(ram16sdp_inst_186_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1028 (
  .O(mux_o_1028),
  .I0(ram16sdp_inst_194_dout[8]),
  .I1(ram16sdp_inst_202_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1029 (
  .O(mux_o_1029),
  .I0(ram16sdp_inst_210_dout[8]),
  .I1(ram16sdp_inst_218_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1030 (
  .O(mux_o_1030),
  .I0(ram16sdp_inst_226_dout[8]),
  .I1(ram16sdp_inst_234_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1031 (
  .O(mux_o_1031),
  .I0(ram16sdp_inst_242_dout[8]),
  .I1(ram16sdp_inst_250_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1032 (
  .O(mux_o_1032),
  .I0(ram16sdp_inst_258_dout[8]),
  .I1(ram16sdp_inst_266_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1033 (
  .O(mux_o_1033),
  .I0(ram16sdp_inst_274_dout[8]),
  .I1(ram16sdp_inst_282_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1034 (
  .O(mux_o_1034),
  .I0(ram16sdp_inst_290_dout[8]),
  .I1(ram16sdp_inst_298_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1035 (
  .O(mux_o_1035),
  .I0(ram16sdp_inst_306_dout[8]),
  .I1(ram16sdp_inst_314_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1036 (
  .O(mux_o_1036),
  .I0(ram16sdp_inst_322_dout[8]),
  .I1(ram16sdp_inst_330_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1037 (
  .O(mux_o_1037),
  .I0(ram16sdp_inst_338_dout[8]),
  .I1(ram16sdp_inst_346_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1038 (
  .O(mux_o_1038),
  .I0(ram16sdp_inst_354_dout[8]),
  .I1(ram16sdp_inst_362_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1039 (
  .O(mux_o_1039),
  .I0(ram16sdp_inst_370_dout[8]),
  .I1(ram16sdp_inst_378_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1040 (
  .O(mux_o_1040),
  .I0(ram16sdp_inst_386_dout[8]),
  .I1(ram16sdp_inst_394_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1041 (
  .O(mux_o_1041),
  .I0(ram16sdp_inst_402_dout[8]),
  .I1(ram16sdp_inst_410_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1042 (
  .O(mux_o_1042),
  .I0(ram16sdp_inst_418_dout[8]),
  .I1(ram16sdp_inst_426_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1043 (
  .O(mux_o_1043),
  .I0(ram16sdp_inst_434_dout[8]),
  .I1(ram16sdp_inst_442_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1044 (
  .O(mux_o_1044),
  .I0(ram16sdp_inst_450_dout[8]),
  .I1(ram16sdp_inst_458_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1045 (
  .O(mux_o_1045),
  .I0(ram16sdp_inst_466_dout[8]),
  .I1(ram16sdp_inst_474_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1046 (
  .O(mux_o_1046),
  .I0(ram16sdp_inst_482_dout[8]),
  .I1(ram16sdp_inst_490_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1047 (
  .O(mux_o_1047),
  .I0(ram16sdp_inst_498_dout[8]),
  .I1(ram16sdp_inst_506_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1048 (
  .O(mux_o_1048),
  .I0(ram16sdp_inst_514_dout[8]),
  .I1(ram16sdp_inst_522_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1049 (
  .O(mux_o_1049),
  .I0(ram16sdp_inst_530_dout[8]),
  .I1(ram16sdp_inst_538_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1050 (
  .O(mux_o_1050),
  .I0(ram16sdp_inst_546_dout[8]),
  .I1(ram16sdp_inst_554_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1051 (
  .O(mux_o_1051),
  .I0(ram16sdp_inst_562_dout[8]),
  .I1(ram16sdp_inst_570_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1052 (
  .O(mux_o_1052),
  .I0(ram16sdp_inst_578_dout[8]),
  .I1(ram16sdp_inst_586_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1053 (
  .O(mux_o_1053),
  .I0(ram16sdp_inst_594_dout[8]),
  .I1(ram16sdp_inst_602_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1054 (
  .O(mux_o_1054),
  .I0(ram16sdp_inst_610_dout[8]),
  .I1(ram16sdp_inst_618_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1055 (
  .O(mux_o_1055),
  .I0(ram16sdp_inst_626_dout[8]),
  .I1(ram16sdp_inst_634_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1056 (
  .O(mux_o_1056),
  .I0(ram16sdp_inst_642_dout[8]),
  .I1(ram16sdp_inst_650_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1057 (
  .O(mux_o_1057),
  .I0(ram16sdp_inst_658_dout[8]),
  .I1(ram16sdp_inst_666_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1058 (
  .O(mux_o_1058),
  .I0(ram16sdp_inst_674_dout[8]),
  .I1(ram16sdp_inst_682_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1059 (
  .O(mux_o_1059),
  .I0(ram16sdp_inst_690_dout[8]),
  .I1(ram16sdp_inst_698_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1060 (
  .O(mux_o_1060),
  .I0(ram16sdp_inst_706_dout[8]),
  .I1(ram16sdp_inst_714_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1061 (
  .O(mux_o_1061),
  .I0(ram16sdp_inst_722_dout[8]),
  .I1(ram16sdp_inst_730_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1062 (
  .O(mux_o_1062),
  .I0(ram16sdp_inst_738_dout[8]),
  .I1(ram16sdp_inst_746_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1063 (
  .O(mux_o_1063),
  .I0(ram16sdp_inst_754_dout[8]),
  .I1(ram16sdp_inst_762_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1064 (
  .O(mux_o_1064),
  .I0(ram16sdp_inst_770_dout[8]),
  .I1(ram16sdp_inst_778_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1065 (
  .O(mux_o_1065),
  .I0(ram16sdp_inst_786_dout[8]),
  .I1(ram16sdp_inst_794_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1066 (
  .O(mux_o_1066),
  .I0(ram16sdp_inst_802_dout[8]),
  .I1(ram16sdp_inst_810_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1067 (
  .O(mux_o_1067),
  .I0(ram16sdp_inst_818_dout[8]),
  .I1(ram16sdp_inst_826_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1068 (
  .O(mux_o_1068),
  .I0(ram16sdp_inst_834_dout[8]),
  .I1(ram16sdp_inst_842_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1069 (
  .O(mux_o_1069),
  .I0(ram16sdp_inst_850_dout[8]),
  .I1(ram16sdp_inst_858_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1070 (
  .O(mux_o_1070),
  .I0(ram16sdp_inst_866_dout[8]),
  .I1(ram16sdp_inst_874_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1071 (
  .O(mux_o_1071),
  .I0(ram16sdp_inst_882_dout[8]),
  .I1(ram16sdp_inst_890_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1072 (
  .O(mux_o_1072),
  .I0(ram16sdp_inst_898_dout[8]),
  .I1(ram16sdp_inst_906_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1073 (
  .O(mux_o_1073),
  .I0(ram16sdp_inst_914_dout[8]),
  .I1(ram16sdp_inst_922_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1074 (
  .O(mux_o_1074),
  .I0(ram16sdp_inst_930_dout[8]),
  .I1(ram16sdp_inst_938_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1075 (
  .O(mux_o_1075),
  .I0(ram16sdp_inst_946_dout[8]),
  .I1(ram16sdp_inst_954_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1076 (
  .O(mux_o_1076),
  .I0(ram16sdp_inst_962_dout[8]),
  .I1(ram16sdp_inst_970_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1077 (
  .O(mux_o_1077),
  .I0(ram16sdp_inst_978_dout[8]),
  .I1(ram16sdp_inst_986_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1078 (
  .O(mux_o_1078),
  .I0(ram16sdp_inst_994_dout[8]),
  .I1(ram16sdp_inst_1002_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1079 (
  .O(mux_o_1079),
  .I0(ram16sdp_inst_1010_dout[8]),
  .I1(ram16sdp_inst_1018_dout[8]),
  .S0(rad[4])
);
MUX2 mux_inst_1080 (
  .O(mux_o_1080),
  .I0(mux_o_1016),
  .I1(mux_o_1017),
  .S0(rad[5])
);
MUX2 mux_inst_1081 (
  .O(mux_o_1081),
  .I0(mux_o_1018),
  .I1(mux_o_1019),
  .S0(rad[5])
);
MUX2 mux_inst_1082 (
  .O(mux_o_1082),
  .I0(mux_o_1020),
  .I1(mux_o_1021),
  .S0(rad[5])
);
MUX2 mux_inst_1083 (
  .O(mux_o_1083),
  .I0(mux_o_1022),
  .I1(mux_o_1023),
  .S0(rad[5])
);
MUX2 mux_inst_1084 (
  .O(mux_o_1084),
  .I0(mux_o_1024),
  .I1(mux_o_1025),
  .S0(rad[5])
);
MUX2 mux_inst_1085 (
  .O(mux_o_1085),
  .I0(mux_o_1026),
  .I1(mux_o_1027),
  .S0(rad[5])
);
MUX2 mux_inst_1086 (
  .O(mux_o_1086),
  .I0(mux_o_1028),
  .I1(mux_o_1029),
  .S0(rad[5])
);
MUX2 mux_inst_1087 (
  .O(mux_o_1087),
  .I0(mux_o_1030),
  .I1(mux_o_1031),
  .S0(rad[5])
);
MUX2 mux_inst_1088 (
  .O(mux_o_1088),
  .I0(mux_o_1032),
  .I1(mux_o_1033),
  .S0(rad[5])
);
MUX2 mux_inst_1089 (
  .O(mux_o_1089),
  .I0(mux_o_1034),
  .I1(mux_o_1035),
  .S0(rad[5])
);
MUX2 mux_inst_1090 (
  .O(mux_o_1090),
  .I0(mux_o_1036),
  .I1(mux_o_1037),
  .S0(rad[5])
);
MUX2 mux_inst_1091 (
  .O(mux_o_1091),
  .I0(mux_o_1038),
  .I1(mux_o_1039),
  .S0(rad[5])
);
MUX2 mux_inst_1092 (
  .O(mux_o_1092),
  .I0(mux_o_1040),
  .I1(mux_o_1041),
  .S0(rad[5])
);
MUX2 mux_inst_1093 (
  .O(mux_o_1093),
  .I0(mux_o_1042),
  .I1(mux_o_1043),
  .S0(rad[5])
);
MUX2 mux_inst_1094 (
  .O(mux_o_1094),
  .I0(mux_o_1044),
  .I1(mux_o_1045),
  .S0(rad[5])
);
MUX2 mux_inst_1095 (
  .O(mux_o_1095),
  .I0(mux_o_1046),
  .I1(mux_o_1047),
  .S0(rad[5])
);
MUX2 mux_inst_1096 (
  .O(mux_o_1096),
  .I0(mux_o_1048),
  .I1(mux_o_1049),
  .S0(rad[5])
);
MUX2 mux_inst_1097 (
  .O(mux_o_1097),
  .I0(mux_o_1050),
  .I1(mux_o_1051),
  .S0(rad[5])
);
MUX2 mux_inst_1098 (
  .O(mux_o_1098),
  .I0(mux_o_1052),
  .I1(mux_o_1053),
  .S0(rad[5])
);
MUX2 mux_inst_1099 (
  .O(mux_o_1099),
  .I0(mux_o_1054),
  .I1(mux_o_1055),
  .S0(rad[5])
);
MUX2 mux_inst_1100 (
  .O(mux_o_1100),
  .I0(mux_o_1056),
  .I1(mux_o_1057),
  .S0(rad[5])
);
MUX2 mux_inst_1101 (
  .O(mux_o_1101),
  .I0(mux_o_1058),
  .I1(mux_o_1059),
  .S0(rad[5])
);
MUX2 mux_inst_1102 (
  .O(mux_o_1102),
  .I0(mux_o_1060),
  .I1(mux_o_1061),
  .S0(rad[5])
);
MUX2 mux_inst_1103 (
  .O(mux_o_1103),
  .I0(mux_o_1062),
  .I1(mux_o_1063),
  .S0(rad[5])
);
MUX2 mux_inst_1104 (
  .O(mux_o_1104),
  .I0(mux_o_1064),
  .I1(mux_o_1065),
  .S0(rad[5])
);
MUX2 mux_inst_1105 (
  .O(mux_o_1105),
  .I0(mux_o_1066),
  .I1(mux_o_1067),
  .S0(rad[5])
);
MUX2 mux_inst_1106 (
  .O(mux_o_1106),
  .I0(mux_o_1068),
  .I1(mux_o_1069),
  .S0(rad[5])
);
MUX2 mux_inst_1107 (
  .O(mux_o_1107),
  .I0(mux_o_1070),
  .I1(mux_o_1071),
  .S0(rad[5])
);
MUX2 mux_inst_1108 (
  .O(mux_o_1108),
  .I0(mux_o_1072),
  .I1(mux_o_1073),
  .S0(rad[5])
);
MUX2 mux_inst_1109 (
  .O(mux_o_1109),
  .I0(mux_o_1074),
  .I1(mux_o_1075),
  .S0(rad[5])
);
MUX2 mux_inst_1110 (
  .O(mux_o_1110),
  .I0(mux_o_1076),
  .I1(mux_o_1077),
  .S0(rad[5])
);
MUX2 mux_inst_1111 (
  .O(mux_o_1111),
  .I0(mux_o_1078),
  .I1(mux_o_1079),
  .S0(rad[5])
);
MUX2 mux_inst_1112 (
  .O(mux_o_1112),
  .I0(mux_o_1080),
  .I1(mux_o_1081),
  .S0(rad[6])
);
MUX2 mux_inst_1113 (
  .O(mux_o_1113),
  .I0(mux_o_1082),
  .I1(mux_o_1083),
  .S0(rad[6])
);
MUX2 mux_inst_1114 (
  .O(mux_o_1114),
  .I0(mux_o_1084),
  .I1(mux_o_1085),
  .S0(rad[6])
);
MUX2 mux_inst_1115 (
  .O(mux_o_1115),
  .I0(mux_o_1086),
  .I1(mux_o_1087),
  .S0(rad[6])
);
MUX2 mux_inst_1116 (
  .O(mux_o_1116),
  .I0(mux_o_1088),
  .I1(mux_o_1089),
  .S0(rad[6])
);
MUX2 mux_inst_1117 (
  .O(mux_o_1117),
  .I0(mux_o_1090),
  .I1(mux_o_1091),
  .S0(rad[6])
);
MUX2 mux_inst_1118 (
  .O(mux_o_1118),
  .I0(mux_o_1092),
  .I1(mux_o_1093),
  .S0(rad[6])
);
MUX2 mux_inst_1119 (
  .O(mux_o_1119),
  .I0(mux_o_1094),
  .I1(mux_o_1095),
  .S0(rad[6])
);
MUX2 mux_inst_1120 (
  .O(mux_o_1120),
  .I0(mux_o_1096),
  .I1(mux_o_1097),
  .S0(rad[6])
);
MUX2 mux_inst_1121 (
  .O(mux_o_1121),
  .I0(mux_o_1098),
  .I1(mux_o_1099),
  .S0(rad[6])
);
MUX2 mux_inst_1122 (
  .O(mux_o_1122),
  .I0(mux_o_1100),
  .I1(mux_o_1101),
  .S0(rad[6])
);
MUX2 mux_inst_1123 (
  .O(mux_o_1123),
  .I0(mux_o_1102),
  .I1(mux_o_1103),
  .S0(rad[6])
);
MUX2 mux_inst_1124 (
  .O(mux_o_1124),
  .I0(mux_o_1104),
  .I1(mux_o_1105),
  .S0(rad[6])
);
MUX2 mux_inst_1125 (
  .O(mux_o_1125),
  .I0(mux_o_1106),
  .I1(mux_o_1107),
  .S0(rad[6])
);
MUX2 mux_inst_1126 (
  .O(mux_o_1126),
  .I0(mux_o_1108),
  .I1(mux_o_1109),
  .S0(rad[6])
);
MUX2 mux_inst_1127 (
  .O(mux_o_1127),
  .I0(mux_o_1110),
  .I1(mux_o_1111),
  .S0(rad[6])
);
MUX2 mux_inst_1128 (
  .O(mux_o_1128),
  .I0(mux_o_1112),
  .I1(mux_o_1113),
  .S0(rad[7])
);
MUX2 mux_inst_1129 (
  .O(mux_o_1129),
  .I0(mux_o_1114),
  .I1(mux_o_1115),
  .S0(rad[7])
);
MUX2 mux_inst_1130 (
  .O(mux_o_1130),
  .I0(mux_o_1116),
  .I1(mux_o_1117),
  .S0(rad[7])
);
MUX2 mux_inst_1131 (
  .O(mux_o_1131),
  .I0(mux_o_1118),
  .I1(mux_o_1119),
  .S0(rad[7])
);
MUX2 mux_inst_1132 (
  .O(mux_o_1132),
  .I0(mux_o_1120),
  .I1(mux_o_1121),
  .S0(rad[7])
);
MUX2 mux_inst_1133 (
  .O(mux_o_1133),
  .I0(mux_o_1122),
  .I1(mux_o_1123),
  .S0(rad[7])
);
MUX2 mux_inst_1134 (
  .O(mux_o_1134),
  .I0(mux_o_1124),
  .I1(mux_o_1125),
  .S0(rad[7])
);
MUX2 mux_inst_1135 (
  .O(mux_o_1135),
  .I0(mux_o_1126),
  .I1(mux_o_1127),
  .S0(rad[7])
);
MUX2 mux_inst_1136 (
  .O(mux_o_1136),
  .I0(mux_o_1128),
  .I1(mux_o_1129),
  .S0(rad[8])
);
MUX2 mux_inst_1137 (
  .O(mux_o_1137),
  .I0(mux_o_1130),
  .I1(mux_o_1131),
  .S0(rad[8])
);
MUX2 mux_inst_1138 (
  .O(mux_o_1138),
  .I0(mux_o_1132),
  .I1(mux_o_1133),
  .S0(rad[8])
);
MUX2 mux_inst_1139 (
  .O(mux_o_1139),
  .I0(mux_o_1134),
  .I1(mux_o_1135),
  .S0(rad[8])
);
MUX2 mux_inst_1140 (
  .O(mux_o_1140),
  .I0(mux_o_1136),
  .I1(mux_o_1137),
  .S0(rad[9])
);
MUX2 mux_inst_1141 (
  .O(mux_o_1141),
  .I0(mux_o_1138),
  .I1(mux_o_1139),
  .S0(rad[9])
);
MUX2 mux_inst_1142 (
  .O(dout[8]),
  .I0(mux_o_1140),
  .I1(mux_o_1141),
  .S0(rad[10])
);
MUX2 mux_inst_1143 (
  .O(mux_o_1143),
  .I0(ram16sdp_inst_2_dout[9]),
  .I1(ram16sdp_inst_10_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1144 (
  .O(mux_o_1144),
  .I0(ram16sdp_inst_18_dout[9]),
  .I1(ram16sdp_inst_26_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1145 (
  .O(mux_o_1145),
  .I0(ram16sdp_inst_34_dout[9]),
  .I1(ram16sdp_inst_42_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1146 (
  .O(mux_o_1146),
  .I0(ram16sdp_inst_50_dout[9]),
  .I1(ram16sdp_inst_58_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1147 (
  .O(mux_o_1147),
  .I0(ram16sdp_inst_66_dout[9]),
  .I1(ram16sdp_inst_74_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1148 (
  .O(mux_o_1148),
  .I0(ram16sdp_inst_82_dout[9]),
  .I1(ram16sdp_inst_90_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1149 (
  .O(mux_o_1149),
  .I0(ram16sdp_inst_98_dout[9]),
  .I1(ram16sdp_inst_106_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1150 (
  .O(mux_o_1150),
  .I0(ram16sdp_inst_114_dout[9]),
  .I1(ram16sdp_inst_122_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1151 (
  .O(mux_o_1151),
  .I0(ram16sdp_inst_130_dout[9]),
  .I1(ram16sdp_inst_138_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1152 (
  .O(mux_o_1152),
  .I0(ram16sdp_inst_146_dout[9]),
  .I1(ram16sdp_inst_154_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1153 (
  .O(mux_o_1153),
  .I0(ram16sdp_inst_162_dout[9]),
  .I1(ram16sdp_inst_170_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1154 (
  .O(mux_o_1154),
  .I0(ram16sdp_inst_178_dout[9]),
  .I1(ram16sdp_inst_186_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1155 (
  .O(mux_o_1155),
  .I0(ram16sdp_inst_194_dout[9]),
  .I1(ram16sdp_inst_202_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1156 (
  .O(mux_o_1156),
  .I0(ram16sdp_inst_210_dout[9]),
  .I1(ram16sdp_inst_218_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1157 (
  .O(mux_o_1157),
  .I0(ram16sdp_inst_226_dout[9]),
  .I1(ram16sdp_inst_234_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1158 (
  .O(mux_o_1158),
  .I0(ram16sdp_inst_242_dout[9]),
  .I1(ram16sdp_inst_250_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1159 (
  .O(mux_o_1159),
  .I0(ram16sdp_inst_258_dout[9]),
  .I1(ram16sdp_inst_266_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1160 (
  .O(mux_o_1160),
  .I0(ram16sdp_inst_274_dout[9]),
  .I1(ram16sdp_inst_282_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1161 (
  .O(mux_o_1161),
  .I0(ram16sdp_inst_290_dout[9]),
  .I1(ram16sdp_inst_298_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1162 (
  .O(mux_o_1162),
  .I0(ram16sdp_inst_306_dout[9]),
  .I1(ram16sdp_inst_314_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1163 (
  .O(mux_o_1163),
  .I0(ram16sdp_inst_322_dout[9]),
  .I1(ram16sdp_inst_330_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1164 (
  .O(mux_o_1164),
  .I0(ram16sdp_inst_338_dout[9]),
  .I1(ram16sdp_inst_346_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1165 (
  .O(mux_o_1165),
  .I0(ram16sdp_inst_354_dout[9]),
  .I1(ram16sdp_inst_362_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1166 (
  .O(mux_o_1166),
  .I0(ram16sdp_inst_370_dout[9]),
  .I1(ram16sdp_inst_378_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1167 (
  .O(mux_o_1167),
  .I0(ram16sdp_inst_386_dout[9]),
  .I1(ram16sdp_inst_394_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1168 (
  .O(mux_o_1168),
  .I0(ram16sdp_inst_402_dout[9]),
  .I1(ram16sdp_inst_410_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1169 (
  .O(mux_o_1169),
  .I0(ram16sdp_inst_418_dout[9]),
  .I1(ram16sdp_inst_426_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1170 (
  .O(mux_o_1170),
  .I0(ram16sdp_inst_434_dout[9]),
  .I1(ram16sdp_inst_442_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1171 (
  .O(mux_o_1171),
  .I0(ram16sdp_inst_450_dout[9]),
  .I1(ram16sdp_inst_458_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1172 (
  .O(mux_o_1172),
  .I0(ram16sdp_inst_466_dout[9]),
  .I1(ram16sdp_inst_474_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1173 (
  .O(mux_o_1173),
  .I0(ram16sdp_inst_482_dout[9]),
  .I1(ram16sdp_inst_490_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1174 (
  .O(mux_o_1174),
  .I0(ram16sdp_inst_498_dout[9]),
  .I1(ram16sdp_inst_506_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1175 (
  .O(mux_o_1175),
  .I0(ram16sdp_inst_514_dout[9]),
  .I1(ram16sdp_inst_522_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1176 (
  .O(mux_o_1176),
  .I0(ram16sdp_inst_530_dout[9]),
  .I1(ram16sdp_inst_538_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1177 (
  .O(mux_o_1177),
  .I0(ram16sdp_inst_546_dout[9]),
  .I1(ram16sdp_inst_554_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1178 (
  .O(mux_o_1178),
  .I0(ram16sdp_inst_562_dout[9]),
  .I1(ram16sdp_inst_570_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1179 (
  .O(mux_o_1179),
  .I0(ram16sdp_inst_578_dout[9]),
  .I1(ram16sdp_inst_586_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1180 (
  .O(mux_o_1180),
  .I0(ram16sdp_inst_594_dout[9]),
  .I1(ram16sdp_inst_602_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1181 (
  .O(mux_o_1181),
  .I0(ram16sdp_inst_610_dout[9]),
  .I1(ram16sdp_inst_618_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1182 (
  .O(mux_o_1182),
  .I0(ram16sdp_inst_626_dout[9]),
  .I1(ram16sdp_inst_634_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1183 (
  .O(mux_o_1183),
  .I0(ram16sdp_inst_642_dout[9]),
  .I1(ram16sdp_inst_650_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1184 (
  .O(mux_o_1184),
  .I0(ram16sdp_inst_658_dout[9]),
  .I1(ram16sdp_inst_666_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1185 (
  .O(mux_o_1185),
  .I0(ram16sdp_inst_674_dout[9]),
  .I1(ram16sdp_inst_682_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1186 (
  .O(mux_o_1186),
  .I0(ram16sdp_inst_690_dout[9]),
  .I1(ram16sdp_inst_698_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1187 (
  .O(mux_o_1187),
  .I0(ram16sdp_inst_706_dout[9]),
  .I1(ram16sdp_inst_714_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1188 (
  .O(mux_o_1188),
  .I0(ram16sdp_inst_722_dout[9]),
  .I1(ram16sdp_inst_730_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1189 (
  .O(mux_o_1189),
  .I0(ram16sdp_inst_738_dout[9]),
  .I1(ram16sdp_inst_746_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1190 (
  .O(mux_o_1190),
  .I0(ram16sdp_inst_754_dout[9]),
  .I1(ram16sdp_inst_762_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1191 (
  .O(mux_o_1191),
  .I0(ram16sdp_inst_770_dout[9]),
  .I1(ram16sdp_inst_778_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1192 (
  .O(mux_o_1192),
  .I0(ram16sdp_inst_786_dout[9]),
  .I1(ram16sdp_inst_794_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1193 (
  .O(mux_o_1193),
  .I0(ram16sdp_inst_802_dout[9]),
  .I1(ram16sdp_inst_810_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1194 (
  .O(mux_o_1194),
  .I0(ram16sdp_inst_818_dout[9]),
  .I1(ram16sdp_inst_826_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1195 (
  .O(mux_o_1195),
  .I0(ram16sdp_inst_834_dout[9]),
  .I1(ram16sdp_inst_842_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1196 (
  .O(mux_o_1196),
  .I0(ram16sdp_inst_850_dout[9]),
  .I1(ram16sdp_inst_858_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1197 (
  .O(mux_o_1197),
  .I0(ram16sdp_inst_866_dout[9]),
  .I1(ram16sdp_inst_874_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1198 (
  .O(mux_o_1198),
  .I0(ram16sdp_inst_882_dout[9]),
  .I1(ram16sdp_inst_890_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1199 (
  .O(mux_o_1199),
  .I0(ram16sdp_inst_898_dout[9]),
  .I1(ram16sdp_inst_906_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1200 (
  .O(mux_o_1200),
  .I0(ram16sdp_inst_914_dout[9]),
  .I1(ram16sdp_inst_922_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1201 (
  .O(mux_o_1201),
  .I0(ram16sdp_inst_930_dout[9]),
  .I1(ram16sdp_inst_938_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1202 (
  .O(mux_o_1202),
  .I0(ram16sdp_inst_946_dout[9]),
  .I1(ram16sdp_inst_954_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1203 (
  .O(mux_o_1203),
  .I0(ram16sdp_inst_962_dout[9]),
  .I1(ram16sdp_inst_970_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1204 (
  .O(mux_o_1204),
  .I0(ram16sdp_inst_978_dout[9]),
  .I1(ram16sdp_inst_986_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1205 (
  .O(mux_o_1205),
  .I0(ram16sdp_inst_994_dout[9]),
  .I1(ram16sdp_inst_1002_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1206 (
  .O(mux_o_1206),
  .I0(ram16sdp_inst_1010_dout[9]),
  .I1(ram16sdp_inst_1018_dout[9]),
  .S0(rad[4])
);
MUX2 mux_inst_1207 (
  .O(mux_o_1207),
  .I0(mux_o_1143),
  .I1(mux_o_1144),
  .S0(rad[5])
);
MUX2 mux_inst_1208 (
  .O(mux_o_1208),
  .I0(mux_o_1145),
  .I1(mux_o_1146),
  .S0(rad[5])
);
MUX2 mux_inst_1209 (
  .O(mux_o_1209),
  .I0(mux_o_1147),
  .I1(mux_o_1148),
  .S0(rad[5])
);
MUX2 mux_inst_1210 (
  .O(mux_o_1210),
  .I0(mux_o_1149),
  .I1(mux_o_1150),
  .S0(rad[5])
);
MUX2 mux_inst_1211 (
  .O(mux_o_1211),
  .I0(mux_o_1151),
  .I1(mux_o_1152),
  .S0(rad[5])
);
MUX2 mux_inst_1212 (
  .O(mux_o_1212),
  .I0(mux_o_1153),
  .I1(mux_o_1154),
  .S0(rad[5])
);
MUX2 mux_inst_1213 (
  .O(mux_o_1213),
  .I0(mux_o_1155),
  .I1(mux_o_1156),
  .S0(rad[5])
);
MUX2 mux_inst_1214 (
  .O(mux_o_1214),
  .I0(mux_o_1157),
  .I1(mux_o_1158),
  .S0(rad[5])
);
MUX2 mux_inst_1215 (
  .O(mux_o_1215),
  .I0(mux_o_1159),
  .I1(mux_o_1160),
  .S0(rad[5])
);
MUX2 mux_inst_1216 (
  .O(mux_o_1216),
  .I0(mux_o_1161),
  .I1(mux_o_1162),
  .S0(rad[5])
);
MUX2 mux_inst_1217 (
  .O(mux_o_1217),
  .I0(mux_o_1163),
  .I1(mux_o_1164),
  .S0(rad[5])
);
MUX2 mux_inst_1218 (
  .O(mux_o_1218),
  .I0(mux_o_1165),
  .I1(mux_o_1166),
  .S0(rad[5])
);
MUX2 mux_inst_1219 (
  .O(mux_o_1219),
  .I0(mux_o_1167),
  .I1(mux_o_1168),
  .S0(rad[5])
);
MUX2 mux_inst_1220 (
  .O(mux_o_1220),
  .I0(mux_o_1169),
  .I1(mux_o_1170),
  .S0(rad[5])
);
MUX2 mux_inst_1221 (
  .O(mux_o_1221),
  .I0(mux_o_1171),
  .I1(mux_o_1172),
  .S0(rad[5])
);
MUX2 mux_inst_1222 (
  .O(mux_o_1222),
  .I0(mux_o_1173),
  .I1(mux_o_1174),
  .S0(rad[5])
);
MUX2 mux_inst_1223 (
  .O(mux_o_1223),
  .I0(mux_o_1175),
  .I1(mux_o_1176),
  .S0(rad[5])
);
MUX2 mux_inst_1224 (
  .O(mux_o_1224),
  .I0(mux_o_1177),
  .I1(mux_o_1178),
  .S0(rad[5])
);
MUX2 mux_inst_1225 (
  .O(mux_o_1225),
  .I0(mux_o_1179),
  .I1(mux_o_1180),
  .S0(rad[5])
);
MUX2 mux_inst_1226 (
  .O(mux_o_1226),
  .I0(mux_o_1181),
  .I1(mux_o_1182),
  .S0(rad[5])
);
MUX2 mux_inst_1227 (
  .O(mux_o_1227),
  .I0(mux_o_1183),
  .I1(mux_o_1184),
  .S0(rad[5])
);
MUX2 mux_inst_1228 (
  .O(mux_o_1228),
  .I0(mux_o_1185),
  .I1(mux_o_1186),
  .S0(rad[5])
);
MUX2 mux_inst_1229 (
  .O(mux_o_1229),
  .I0(mux_o_1187),
  .I1(mux_o_1188),
  .S0(rad[5])
);
MUX2 mux_inst_1230 (
  .O(mux_o_1230),
  .I0(mux_o_1189),
  .I1(mux_o_1190),
  .S0(rad[5])
);
MUX2 mux_inst_1231 (
  .O(mux_o_1231),
  .I0(mux_o_1191),
  .I1(mux_o_1192),
  .S0(rad[5])
);
MUX2 mux_inst_1232 (
  .O(mux_o_1232),
  .I0(mux_o_1193),
  .I1(mux_o_1194),
  .S0(rad[5])
);
MUX2 mux_inst_1233 (
  .O(mux_o_1233),
  .I0(mux_o_1195),
  .I1(mux_o_1196),
  .S0(rad[5])
);
MUX2 mux_inst_1234 (
  .O(mux_o_1234),
  .I0(mux_o_1197),
  .I1(mux_o_1198),
  .S0(rad[5])
);
MUX2 mux_inst_1235 (
  .O(mux_o_1235),
  .I0(mux_o_1199),
  .I1(mux_o_1200),
  .S0(rad[5])
);
MUX2 mux_inst_1236 (
  .O(mux_o_1236),
  .I0(mux_o_1201),
  .I1(mux_o_1202),
  .S0(rad[5])
);
MUX2 mux_inst_1237 (
  .O(mux_o_1237),
  .I0(mux_o_1203),
  .I1(mux_o_1204),
  .S0(rad[5])
);
MUX2 mux_inst_1238 (
  .O(mux_o_1238),
  .I0(mux_o_1205),
  .I1(mux_o_1206),
  .S0(rad[5])
);
MUX2 mux_inst_1239 (
  .O(mux_o_1239),
  .I0(mux_o_1207),
  .I1(mux_o_1208),
  .S0(rad[6])
);
MUX2 mux_inst_1240 (
  .O(mux_o_1240),
  .I0(mux_o_1209),
  .I1(mux_o_1210),
  .S0(rad[6])
);
MUX2 mux_inst_1241 (
  .O(mux_o_1241),
  .I0(mux_o_1211),
  .I1(mux_o_1212),
  .S0(rad[6])
);
MUX2 mux_inst_1242 (
  .O(mux_o_1242),
  .I0(mux_o_1213),
  .I1(mux_o_1214),
  .S0(rad[6])
);
MUX2 mux_inst_1243 (
  .O(mux_o_1243),
  .I0(mux_o_1215),
  .I1(mux_o_1216),
  .S0(rad[6])
);
MUX2 mux_inst_1244 (
  .O(mux_o_1244),
  .I0(mux_o_1217),
  .I1(mux_o_1218),
  .S0(rad[6])
);
MUX2 mux_inst_1245 (
  .O(mux_o_1245),
  .I0(mux_o_1219),
  .I1(mux_o_1220),
  .S0(rad[6])
);
MUX2 mux_inst_1246 (
  .O(mux_o_1246),
  .I0(mux_o_1221),
  .I1(mux_o_1222),
  .S0(rad[6])
);
MUX2 mux_inst_1247 (
  .O(mux_o_1247),
  .I0(mux_o_1223),
  .I1(mux_o_1224),
  .S0(rad[6])
);
MUX2 mux_inst_1248 (
  .O(mux_o_1248),
  .I0(mux_o_1225),
  .I1(mux_o_1226),
  .S0(rad[6])
);
MUX2 mux_inst_1249 (
  .O(mux_o_1249),
  .I0(mux_o_1227),
  .I1(mux_o_1228),
  .S0(rad[6])
);
MUX2 mux_inst_1250 (
  .O(mux_o_1250),
  .I0(mux_o_1229),
  .I1(mux_o_1230),
  .S0(rad[6])
);
MUX2 mux_inst_1251 (
  .O(mux_o_1251),
  .I0(mux_o_1231),
  .I1(mux_o_1232),
  .S0(rad[6])
);
MUX2 mux_inst_1252 (
  .O(mux_o_1252),
  .I0(mux_o_1233),
  .I1(mux_o_1234),
  .S0(rad[6])
);
MUX2 mux_inst_1253 (
  .O(mux_o_1253),
  .I0(mux_o_1235),
  .I1(mux_o_1236),
  .S0(rad[6])
);
MUX2 mux_inst_1254 (
  .O(mux_o_1254),
  .I0(mux_o_1237),
  .I1(mux_o_1238),
  .S0(rad[6])
);
MUX2 mux_inst_1255 (
  .O(mux_o_1255),
  .I0(mux_o_1239),
  .I1(mux_o_1240),
  .S0(rad[7])
);
MUX2 mux_inst_1256 (
  .O(mux_o_1256),
  .I0(mux_o_1241),
  .I1(mux_o_1242),
  .S0(rad[7])
);
MUX2 mux_inst_1257 (
  .O(mux_o_1257),
  .I0(mux_o_1243),
  .I1(mux_o_1244),
  .S0(rad[7])
);
MUX2 mux_inst_1258 (
  .O(mux_o_1258),
  .I0(mux_o_1245),
  .I1(mux_o_1246),
  .S0(rad[7])
);
MUX2 mux_inst_1259 (
  .O(mux_o_1259),
  .I0(mux_o_1247),
  .I1(mux_o_1248),
  .S0(rad[7])
);
MUX2 mux_inst_1260 (
  .O(mux_o_1260),
  .I0(mux_o_1249),
  .I1(mux_o_1250),
  .S0(rad[7])
);
MUX2 mux_inst_1261 (
  .O(mux_o_1261),
  .I0(mux_o_1251),
  .I1(mux_o_1252),
  .S0(rad[7])
);
MUX2 mux_inst_1262 (
  .O(mux_o_1262),
  .I0(mux_o_1253),
  .I1(mux_o_1254),
  .S0(rad[7])
);
MUX2 mux_inst_1263 (
  .O(mux_o_1263),
  .I0(mux_o_1255),
  .I1(mux_o_1256),
  .S0(rad[8])
);
MUX2 mux_inst_1264 (
  .O(mux_o_1264),
  .I0(mux_o_1257),
  .I1(mux_o_1258),
  .S0(rad[8])
);
MUX2 mux_inst_1265 (
  .O(mux_o_1265),
  .I0(mux_o_1259),
  .I1(mux_o_1260),
  .S0(rad[8])
);
MUX2 mux_inst_1266 (
  .O(mux_o_1266),
  .I0(mux_o_1261),
  .I1(mux_o_1262),
  .S0(rad[8])
);
MUX2 mux_inst_1267 (
  .O(mux_o_1267),
  .I0(mux_o_1263),
  .I1(mux_o_1264),
  .S0(rad[9])
);
MUX2 mux_inst_1268 (
  .O(mux_o_1268),
  .I0(mux_o_1265),
  .I1(mux_o_1266),
  .S0(rad[9])
);
MUX2 mux_inst_1269 (
  .O(dout[9]),
  .I0(mux_o_1267),
  .I1(mux_o_1268),
  .S0(rad[10])
);
MUX2 mux_inst_1270 (
  .O(mux_o_1270),
  .I0(ram16sdp_inst_2_dout[10]),
  .I1(ram16sdp_inst_10_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1271 (
  .O(mux_o_1271),
  .I0(ram16sdp_inst_18_dout[10]),
  .I1(ram16sdp_inst_26_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1272 (
  .O(mux_o_1272),
  .I0(ram16sdp_inst_34_dout[10]),
  .I1(ram16sdp_inst_42_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1273 (
  .O(mux_o_1273),
  .I0(ram16sdp_inst_50_dout[10]),
  .I1(ram16sdp_inst_58_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1274 (
  .O(mux_o_1274),
  .I0(ram16sdp_inst_66_dout[10]),
  .I1(ram16sdp_inst_74_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1275 (
  .O(mux_o_1275),
  .I0(ram16sdp_inst_82_dout[10]),
  .I1(ram16sdp_inst_90_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1276 (
  .O(mux_o_1276),
  .I0(ram16sdp_inst_98_dout[10]),
  .I1(ram16sdp_inst_106_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1277 (
  .O(mux_o_1277),
  .I0(ram16sdp_inst_114_dout[10]),
  .I1(ram16sdp_inst_122_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1278 (
  .O(mux_o_1278),
  .I0(ram16sdp_inst_130_dout[10]),
  .I1(ram16sdp_inst_138_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1279 (
  .O(mux_o_1279),
  .I0(ram16sdp_inst_146_dout[10]),
  .I1(ram16sdp_inst_154_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1280 (
  .O(mux_o_1280),
  .I0(ram16sdp_inst_162_dout[10]),
  .I1(ram16sdp_inst_170_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1281 (
  .O(mux_o_1281),
  .I0(ram16sdp_inst_178_dout[10]),
  .I1(ram16sdp_inst_186_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1282 (
  .O(mux_o_1282),
  .I0(ram16sdp_inst_194_dout[10]),
  .I1(ram16sdp_inst_202_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1283 (
  .O(mux_o_1283),
  .I0(ram16sdp_inst_210_dout[10]),
  .I1(ram16sdp_inst_218_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1284 (
  .O(mux_o_1284),
  .I0(ram16sdp_inst_226_dout[10]),
  .I1(ram16sdp_inst_234_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1285 (
  .O(mux_o_1285),
  .I0(ram16sdp_inst_242_dout[10]),
  .I1(ram16sdp_inst_250_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1286 (
  .O(mux_o_1286),
  .I0(ram16sdp_inst_258_dout[10]),
  .I1(ram16sdp_inst_266_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1287 (
  .O(mux_o_1287),
  .I0(ram16sdp_inst_274_dout[10]),
  .I1(ram16sdp_inst_282_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1288 (
  .O(mux_o_1288),
  .I0(ram16sdp_inst_290_dout[10]),
  .I1(ram16sdp_inst_298_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1289 (
  .O(mux_o_1289),
  .I0(ram16sdp_inst_306_dout[10]),
  .I1(ram16sdp_inst_314_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1290 (
  .O(mux_o_1290),
  .I0(ram16sdp_inst_322_dout[10]),
  .I1(ram16sdp_inst_330_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1291 (
  .O(mux_o_1291),
  .I0(ram16sdp_inst_338_dout[10]),
  .I1(ram16sdp_inst_346_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1292 (
  .O(mux_o_1292),
  .I0(ram16sdp_inst_354_dout[10]),
  .I1(ram16sdp_inst_362_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1293 (
  .O(mux_o_1293),
  .I0(ram16sdp_inst_370_dout[10]),
  .I1(ram16sdp_inst_378_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1294 (
  .O(mux_o_1294),
  .I0(ram16sdp_inst_386_dout[10]),
  .I1(ram16sdp_inst_394_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1295 (
  .O(mux_o_1295),
  .I0(ram16sdp_inst_402_dout[10]),
  .I1(ram16sdp_inst_410_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1296 (
  .O(mux_o_1296),
  .I0(ram16sdp_inst_418_dout[10]),
  .I1(ram16sdp_inst_426_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1297 (
  .O(mux_o_1297),
  .I0(ram16sdp_inst_434_dout[10]),
  .I1(ram16sdp_inst_442_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1298 (
  .O(mux_o_1298),
  .I0(ram16sdp_inst_450_dout[10]),
  .I1(ram16sdp_inst_458_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1299 (
  .O(mux_o_1299),
  .I0(ram16sdp_inst_466_dout[10]),
  .I1(ram16sdp_inst_474_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1300 (
  .O(mux_o_1300),
  .I0(ram16sdp_inst_482_dout[10]),
  .I1(ram16sdp_inst_490_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1301 (
  .O(mux_o_1301),
  .I0(ram16sdp_inst_498_dout[10]),
  .I1(ram16sdp_inst_506_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1302 (
  .O(mux_o_1302),
  .I0(ram16sdp_inst_514_dout[10]),
  .I1(ram16sdp_inst_522_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1303 (
  .O(mux_o_1303),
  .I0(ram16sdp_inst_530_dout[10]),
  .I1(ram16sdp_inst_538_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1304 (
  .O(mux_o_1304),
  .I0(ram16sdp_inst_546_dout[10]),
  .I1(ram16sdp_inst_554_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1305 (
  .O(mux_o_1305),
  .I0(ram16sdp_inst_562_dout[10]),
  .I1(ram16sdp_inst_570_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1306 (
  .O(mux_o_1306),
  .I0(ram16sdp_inst_578_dout[10]),
  .I1(ram16sdp_inst_586_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1307 (
  .O(mux_o_1307),
  .I0(ram16sdp_inst_594_dout[10]),
  .I1(ram16sdp_inst_602_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1308 (
  .O(mux_o_1308),
  .I0(ram16sdp_inst_610_dout[10]),
  .I1(ram16sdp_inst_618_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1309 (
  .O(mux_o_1309),
  .I0(ram16sdp_inst_626_dout[10]),
  .I1(ram16sdp_inst_634_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1310 (
  .O(mux_o_1310),
  .I0(ram16sdp_inst_642_dout[10]),
  .I1(ram16sdp_inst_650_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1311 (
  .O(mux_o_1311),
  .I0(ram16sdp_inst_658_dout[10]),
  .I1(ram16sdp_inst_666_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1312 (
  .O(mux_o_1312),
  .I0(ram16sdp_inst_674_dout[10]),
  .I1(ram16sdp_inst_682_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1313 (
  .O(mux_o_1313),
  .I0(ram16sdp_inst_690_dout[10]),
  .I1(ram16sdp_inst_698_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1314 (
  .O(mux_o_1314),
  .I0(ram16sdp_inst_706_dout[10]),
  .I1(ram16sdp_inst_714_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1315 (
  .O(mux_o_1315),
  .I0(ram16sdp_inst_722_dout[10]),
  .I1(ram16sdp_inst_730_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1316 (
  .O(mux_o_1316),
  .I0(ram16sdp_inst_738_dout[10]),
  .I1(ram16sdp_inst_746_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1317 (
  .O(mux_o_1317),
  .I0(ram16sdp_inst_754_dout[10]),
  .I1(ram16sdp_inst_762_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1318 (
  .O(mux_o_1318),
  .I0(ram16sdp_inst_770_dout[10]),
  .I1(ram16sdp_inst_778_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1319 (
  .O(mux_o_1319),
  .I0(ram16sdp_inst_786_dout[10]),
  .I1(ram16sdp_inst_794_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1320 (
  .O(mux_o_1320),
  .I0(ram16sdp_inst_802_dout[10]),
  .I1(ram16sdp_inst_810_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1321 (
  .O(mux_o_1321),
  .I0(ram16sdp_inst_818_dout[10]),
  .I1(ram16sdp_inst_826_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1322 (
  .O(mux_o_1322),
  .I0(ram16sdp_inst_834_dout[10]),
  .I1(ram16sdp_inst_842_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1323 (
  .O(mux_o_1323),
  .I0(ram16sdp_inst_850_dout[10]),
  .I1(ram16sdp_inst_858_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1324 (
  .O(mux_o_1324),
  .I0(ram16sdp_inst_866_dout[10]),
  .I1(ram16sdp_inst_874_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1325 (
  .O(mux_o_1325),
  .I0(ram16sdp_inst_882_dout[10]),
  .I1(ram16sdp_inst_890_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1326 (
  .O(mux_o_1326),
  .I0(ram16sdp_inst_898_dout[10]),
  .I1(ram16sdp_inst_906_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1327 (
  .O(mux_o_1327),
  .I0(ram16sdp_inst_914_dout[10]),
  .I1(ram16sdp_inst_922_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1328 (
  .O(mux_o_1328),
  .I0(ram16sdp_inst_930_dout[10]),
  .I1(ram16sdp_inst_938_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1329 (
  .O(mux_o_1329),
  .I0(ram16sdp_inst_946_dout[10]),
  .I1(ram16sdp_inst_954_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1330 (
  .O(mux_o_1330),
  .I0(ram16sdp_inst_962_dout[10]),
  .I1(ram16sdp_inst_970_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1331 (
  .O(mux_o_1331),
  .I0(ram16sdp_inst_978_dout[10]),
  .I1(ram16sdp_inst_986_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1332 (
  .O(mux_o_1332),
  .I0(ram16sdp_inst_994_dout[10]),
  .I1(ram16sdp_inst_1002_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1333 (
  .O(mux_o_1333),
  .I0(ram16sdp_inst_1010_dout[10]),
  .I1(ram16sdp_inst_1018_dout[10]),
  .S0(rad[4])
);
MUX2 mux_inst_1334 (
  .O(mux_o_1334),
  .I0(mux_o_1270),
  .I1(mux_o_1271),
  .S0(rad[5])
);
MUX2 mux_inst_1335 (
  .O(mux_o_1335),
  .I0(mux_o_1272),
  .I1(mux_o_1273),
  .S0(rad[5])
);
MUX2 mux_inst_1336 (
  .O(mux_o_1336),
  .I0(mux_o_1274),
  .I1(mux_o_1275),
  .S0(rad[5])
);
MUX2 mux_inst_1337 (
  .O(mux_o_1337),
  .I0(mux_o_1276),
  .I1(mux_o_1277),
  .S0(rad[5])
);
MUX2 mux_inst_1338 (
  .O(mux_o_1338),
  .I0(mux_o_1278),
  .I1(mux_o_1279),
  .S0(rad[5])
);
MUX2 mux_inst_1339 (
  .O(mux_o_1339),
  .I0(mux_o_1280),
  .I1(mux_o_1281),
  .S0(rad[5])
);
MUX2 mux_inst_1340 (
  .O(mux_o_1340),
  .I0(mux_o_1282),
  .I1(mux_o_1283),
  .S0(rad[5])
);
MUX2 mux_inst_1341 (
  .O(mux_o_1341),
  .I0(mux_o_1284),
  .I1(mux_o_1285),
  .S0(rad[5])
);
MUX2 mux_inst_1342 (
  .O(mux_o_1342),
  .I0(mux_o_1286),
  .I1(mux_o_1287),
  .S0(rad[5])
);
MUX2 mux_inst_1343 (
  .O(mux_o_1343),
  .I0(mux_o_1288),
  .I1(mux_o_1289),
  .S0(rad[5])
);
MUX2 mux_inst_1344 (
  .O(mux_o_1344),
  .I0(mux_o_1290),
  .I1(mux_o_1291),
  .S0(rad[5])
);
MUX2 mux_inst_1345 (
  .O(mux_o_1345),
  .I0(mux_o_1292),
  .I1(mux_o_1293),
  .S0(rad[5])
);
MUX2 mux_inst_1346 (
  .O(mux_o_1346),
  .I0(mux_o_1294),
  .I1(mux_o_1295),
  .S0(rad[5])
);
MUX2 mux_inst_1347 (
  .O(mux_o_1347),
  .I0(mux_o_1296),
  .I1(mux_o_1297),
  .S0(rad[5])
);
MUX2 mux_inst_1348 (
  .O(mux_o_1348),
  .I0(mux_o_1298),
  .I1(mux_o_1299),
  .S0(rad[5])
);
MUX2 mux_inst_1349 (
  .O(mux_o_1349),
  .I0(mux_o_1300),
  .I1(mux_o_1301),
  .S0(rad[5])
);
MUX2 mux_inst_1350 (
  .O(mux_o_1350),
  .I0(mux_o_1302),
  .I1(mux_o_1303),
  .S0(rad[5])
);
MUX2 mux_inst_1351 (
  .O(mux_o_1351),
  .I0(mux_o_1304),
  .I1(mux_o_1305),
  .S0(rad[5])
);
MUX2 mux_inst_1352 (
  .O(mux_o_1352),
  .I0(mux_o_1306),
  .I1(mux_o_1307),
  .S0(rad[5])
);
MUX2 mux_inst_1353 (
  .O(mux_o_1353),
  .I0(mux_o_1308),
  .I1(mux_o_1309),
  .S0(rad[5])
);
MUX2 mux_inst_1354 (
  .O(mux_o_1354),
  .I0(mux_o_1310),
  .I1(mux_o_1311),
  .S0(rad[5])
);
MUX2 mux_inst_1355 (
  .O(mux_o_1355),
  .I0(mux_o_1312),
  .I1(mux_o_1313),
  .S0(rad[5])
);
MUX2 mux_inst_1356 (
  .O(mux_o_1356),
  .I0(mux_o_1314),
  .I1(mux_o_1315),
  .S0(rad[5])
);
MUX2 mux_inst_1357 (
  .O(mux_o_1357),
  .I0(mux_o_1316),
  .I1(mux_o_1317),
  .S0(rad[5])
);
MUX2 mux_inst_1358 (
  .O(mux_o_1358),
  .I0(mux_o_1318),
  .I1(mux_o_1319),
  .S0(rad[5])
);
MUX2 mux_inst_1359 (
  .O(mux_o_1359),
  .I0(mux_o_1320),
  .I1(mux_o_1321),
  .S0(rad[5])
);
MUX2 mux_inst_1360 (
  .O(mux_o_1360),
  .I0(mux_o_1322),
  .I1(mux_o_1323),
  .S0(rad[5])
);
MUX2 mux_inst_1361 (
  .O(mux_o_1361),
  .I0(mux_o_1324),
  .I1(mux_o_1325),
  .S0(rad[5])
);
MUX2 mux_inst_1362 (
  .O(mux_o_1362),
  .I0(mux_o_1326),
  .I1(mux_o_1327),
  .S0(rad[5])
);
MUX2 mux_inst_1363 (
  .O(mux_o_1363),
  .I0(mux_o_1328),
  .I1(mux_o_1329),
  .S0(rad[5])
);
MUX2 mux_inst_1364 (
  .O(mux_o_1364),
  .I0(mux_o_1330),
  .I1(mux_o_1331),
  .S0(rad[5])
);
MUX2 mux_inst_1365 (
  .O(mux_o_1365),
  .I0(mux_o_1332),
  .I1(mux_o_1333),
  .S0(rad[5])
);
MUX2 mux_inst_1366 (
  .O(mux_o_1366),
  .I0(mux_o_1334),
  .I1(mux_o_1335),
  .S0(rad[6])
);
MUX2 mux_inst_1367 (
  .O(mux_o_1367),
  .I0(mux_o_1336),
  .I1(mux_o_1337),
  .S0(rad[6])
);
MUX2 mux_inst_1368 (
  .O(mux_o_1368),
  .I0(mux_o_1338),
  .I1(mux_o_1339),
  .S0(rad[6])
);
MUX2 mux_inst_1369 (
  .O(mux_o_1369),
  .I0(mux_o_1340),
  .I1(mux_o_1341),
  .S0(rad[6])
);
MUX2 mux_inst_1370 (
  .O(mux_o_1370),
  .I0(mux_o_1342),
  .I1(mux_o_1343),
  .S0(rad[6])
);
MUX2 mux_inst_1371 (
  .O(mux_o_1371),
  .I0(mux_o_1344),
  .I1(mux_o_1345),
  .S0(rad[6])
);
MUX2 mux_inst_1372 (
  .O(mux_o_1372),
  .I0(mux_o_1346),
  .I1(mux_o_1347),
  .S0(rad[6])
);
MUX2 mux_inst_1373 (
  .O(mux_o_1373),
  .I0(mux_o_1348),
  .I1(mux_o_1349),
  .S0(rad[6])
);
MUX2 mux_inst_1374 (
  .O(mux_o_1374),
  .I0(mux_o_1350),
  .I1(mux_o_1351),
  .S0(rad[6])
);
MUX2 mux_inst_1375 (
  .O(mux_o_1375),
  .I0(mux_o_1352),
  .I1(mux_o_1353),
  .S0(rad[6])
);
MUX2 mux_inst_1376 (
  .O(mux_o_1376),
  .I0(mux_o_1354),
  .I1(mux_o_1355),
  .S0(rad[6])
);
MUX2 mux_inst_1377 (
  .O(mux_o_1377),
  .I0(mux_o_1356),
  .I1(mux_o_1357),
  .S0(rad[6])
);
MUX2 mux_inst_1378 (
  .O(mux_o_1378),
  .I0(mux_o_1358),
  .I1(mux_o_1359),
  .S0(rad[6])
);
MUX2 mux_inst_1379 (
  .O(mux_o_1379),
  .I0(mux_o_1360),
  .I1(mux_o_1361),
  .S0(rad[6])
);
MUX2 mux_inst_1380 (
  .O(mux_o_1380),
  .I0(mux_o_1362),
  .I1(mux_o_1363),
  .S0(rad[6])
);
MUX2 mux_inst_1381 (
  .O(mux_o_1381),
  .I0(mux_o_1364),
  .I1(mux_o_1365),
  .S0(rad[6])
);
MUX2 mux_inst_1382 (
  .O(mux_o_1382),
  .I0(mux_o_1366),
  .I1(mux_o_1367),
  .S0(rad[7])
);
MUX2 mux_inst_1383 (
  .O(mux_o_1383),
  .I0(mux_o_1368),
  .I1(mux_o_1369),
  .S0(rad[7])
);
MUX2 mux_inst_1384 (
  .O(mux_o_1384),
  .I0(mux_o_1370),
  .I1(mux_o_1371),
  .S0(rad[7])
);
MUX2 mux_inst_1385 (
  .O(mux_o_1385),
  .I0(mux_o_1372),
  .I1(mux_o_1373),
  .S0(rad[7])
);
MUX2 mux_inst_1386 (
  .O(mux_o_1386),
  .I0(mux_o_1374),
  .I1(mux_o_1375),
  .S0(rad[7])
);
MUX2 mux_inst_1387 (
  .O(mux_o_1387),
  .I0(mux_o_1376),
  .I1(mux_o_1377),
  .S0(rad[7])
);
MUX2 mux_inst_1388 (
  .O(mux_o_1388),
  .I0(mux_o_1378),
  .I1(mux_o_1379),
  .S0(rad[7])
);
MUX2 mux_inst_1389 (
  .O(mux_o_1389),
  .I0(mux_o_1380),
  .I1(mux_o_1381),
  .S0(rad[7])
);
MUX2 mux_inst_1390 (
  .O(mux_o_1390),
  .I0(mux_o_1382),
  .I1(mux_o_1383),
  .S0(rad[8])
);
MUX2 mux_inst_1391 (
  .O(mux_o_1391),
  .I0(mux_o_1384),
  .I1(mux_o_1385),
  .S0(rad[8])
);
MUX2 mux_inst_1392 (
  .O(mux_o_1392),
  .I0(mux_o_1386),
  .I1(mux_o_1387),
  .S0(rad[8])
);
MUX2 mux_inst_1393 (
  .O(mux_o_1393),
  .I0(mux_o_1388),
  .I1(mux_o_1389),
  .S0(rad[8])
);
MUX2 mux_inst_1394 (
  .O(mux_o_1394),
  .I0(mux_o_1390),
  .I1(mux_o_1391),
  .S0(rad[9])
);
MUX2 mux_inst_1395 (
  .O(mux_o_1395),
  .I0(mux_o_1392),
  .I1(mux_o_1393),
  .S0(rad[9])
);
MUX2 mux_inst_1396 (
  .O(dout[10]),
  .I0(mux_o_1394),
  .I1(mux_o_1395),
  .S0(rad[10])
);
MUX2 mux_inst_1397 (
  .O(mux_o_1397),
  .I0(ram16sdp_inst_2_dout[11]),
  .I1(ram16sdp_inst_10_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1398 (
  .O(mux_o_1398),
  .I0(ram16sdp_inst_18_dout[11]),
  .I1(ram16sdp_inst_26_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1399 (
  .O(mux_o_1399),
  .I0(ram16sdp_inst_34_dout[11]),
  .I1(ram16sdp_inst_42_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1400 (
  .O(mux_o_1400),
  .I0(ram16sdp_inst_50_dout[11]),
  .I1(ram16sdp_inst_58_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1401 (
  .O(mux_o_1401),
  .I0(ram16sdp_inst_66_dout[11]),
  .I1(ram16sdp_inst_74_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1402 (
  .O(mux_o_1402),
  .I0(ram16sdp_inst_82_dout[11]),
  .I1(ram16sdp_inst_90_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1403 (
  .O(mux_o_1403),
  .I0(ram16sdp_inst_98_dout[11]),
  .I1(ram16sdp_inst_106_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1404 (
  .O(mux_o_1404),
  .I0(ram16sdp_inst_114_dout[11]),
  .I1(ram16sdp_inst_122_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1405 (
  .O(mux_o_1405),
  .I0(ram16sdp_inst_130_dout[11]),
  .I1(ram16sdp_inst_138_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1406 (
  .O(mux_o_1406),
  .I0(ram16sdp_inst_146_dout[11]),
  .I1(ram16sdp_inst_154_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1407 (
  .O(mux_o_1407),
  .I0(ram16sdp_inst_162_dout[11]),
  .I1(ram16sdp_inst_170_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1408 (
  .O(mux_o_1408),
  .I0(ram16sdp_inst_178_dout[11]),
  .I1(ram16sdp_inst_186_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1409 (
  .O(mux_o_1409),
  .I0(ram16sdp_inst_194_dout[11]),
  .I1(ram16sdp_inst_202_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1410 (
  .O(mux_o_1410),
  .I0(ram16sdp_inst_210_dout[11]),
  .I1(ram16sdp_inst_218_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1411 (
  .O(mux_o_1411),
  .I0(ram16sdp_inst_226_dout[11]),
  .I1(ram16sdp_inst_234_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1412 (
  .O(mux_o_1412),
  .I0(ram16sdp_inst_242_dout[11]),
  .I1(ram16sdp_inst_250_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1413 (
  .O(mux_o_1413),
  .I0(ram16sdp_inst_258_dout[11]),
  .I1(ram16sdp_inst_266_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1414 (
  .O(mux_o_1414),
  .I0(ram16sdp_inst_274_dout[11]),
  .I1(ram16sdp_inst_282_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1415 (
  .O(mux_o_1415),
  .I0(ram16sdp_inst_290_dout[11]),
  .I1(ram16sdp_inst_298_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1416 (
  .O(mux_o_1416),
  .I0(ram16sdp_inst_306_dout[11]),
  .I1(ram16sdp_inst_314_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1417 (
  .O(mux_o_1417),
  .I0(ram16sdp_inst_322_dout[11]),
  .I1(ram16sdp_inst_330_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1418 (
  .O(mux_o_1418),
  .I0(ram16sdp_inst_338_dout[11]),
  .I1(ram16sdp_inst_346_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1419 (
  .O(mux_o_1419),
  .I0(ram16sdp_inst_354_dout[11]),
  .I1(ram16sdp_inst_362_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1420 (
  .O(mux_o_1420),
  .I0(ram16sdp_inst_370_dout[11]),
  .I1(ram16sdp_inst_378_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1421 (
  .O(mux_o_1421),
  .I0(ram16sdp_inst_386_dout[11]),
  .I1(ram16sdp_inst_394_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1422 (
  .O(mux_o_1422),
  .I0(ram16sdp_inst_402_dout[11]),
  .I1(ram16sdp_inst_410_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1423 (
  .O(mux_o_1423),
  .I0(ram16sdp_inst_418_dout[11]),
  .I1(ram16sdp_inst_426_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1424 (
  .O(mux_o_1424),
  .I0(ram16sdp_inst_434_dout[11]),
  .I1(ram16sdp_inst_442_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1425 (
  .O(mux_o_1425),
  .I0(ram16sdp_inst_450_dout[11]),
  .I1(ram16sdp_inst_458_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1426 (
  .O(mux_o_1426),
  .I0(ram16sdp_inst_466_dout[11]),
  .I1(ram16sdp_inst_474_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1427 (
  .O(mux_o_1427),
  .I0(ram16sdp_inst_482_dout[11]),
  .I1(ram16sdp_inst_490_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1428 (
  .O(mux_o_1428),
  .I0(ram16sdp_inst_498_dout[11]),
  .I1(ram16sdp_inst_506_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1429 (
  .O(mux_o_1429),
  .I0(ram16sdp_inst_514_dout[11]),
  .I1(ram16sdp_inst_522_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1430 (
  .O(mux_o_1430),
  .I0(ram16sdp_inst_530_dout[11]),
  .I1(ram16sdp_inst_538_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1431 (
  .O(mux_o_1431),
  .I0(ram16sdp_inst_546_dout[11]),
  .I1(ram16sdp_inst_554_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1432 (
  .O(mux_o_1432),
  .I0(ram16sdp_inst_562_dout[11]),
  .I1(ram16sdp_inst_570_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1433 (
  .O(mux_o_1433),
  .I0(ram16sdp_inst_578_dout[11]),
  .I1(ram16sdp_inst_586_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1434 (
  .O(mux_o_1434),
  .I0(ram16sdp_inst_594_dout[11]),
  .I1(ram16sdp_inst_602_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1435 (
  .O(mux_o_1435),
  .I0(ram16sdp_inst_610_dout[11]),
  .I1(ram16sdp_inst_618_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1436 (
  .O(mux_o_1436),
  .I0(ram16sdp_inst_626_dout[11]),
  .I1(ram16sdp_inst_634_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1437 (
  .O(mux_o_1437),
  .I0(ram16sdp_inst_642_dout[11]),
  .I1(ram16sdp_inst_650_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1438 (
  .O(mux_o_1438),
  .I0(ram16sdp_inst_658_dout[11]),
  .I1(ram16sdp_inst_666_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1439 (
  .O(mux_o_1439),
  .I0(ram16sdp_inst_674_dout[11]),
  .I1(ram16sdp_inst_682_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1440 (
  .O(mux_o_1440),
  .I0(ram16sdp_inst_690_dout[11]),
  .I1(ram16sdp_inst_698_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1441 (
  .O(mux_o_1441),
  .I0(ram16sdp_inst_706_dout[11]),
  .I1(ram16sdp_inst_714_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1442 (
  .O(mux_o_1442),
  .I0(ram16sdp_inst_722_dout[11]),
  .I1(ram16sdp_inst_730_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1443 (
  .O(mux_o_1443),
  .I0(ram16sdp_inst_738_dout[11]),
  .I1(ram16sdp_inst_746_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1444 (
  .O(mux_o_1444),
  .I0(ram16sdp_inst_754_dout[11]),
  .I1(ram16sdp_inst_762_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1445 (
  .O(mux_o_1445),
  .I0(ram16sdp_inst_770_dout[11]),
  .I1(ram16sdp_inst_778_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1446 (
  .O(mux_o_1446),
  .I0(ram16sdp_inst_786_dout[11]),
  .I1(ram16sdp_inst_794_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1447 (
  .O(mux_o_1447),
  .I0(ram16sdp_inst_802_dout[11]),
  .I1(ram16sdp_inst_810_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1448 (
  .O(mux_o_1448),
  .I0(ram16sdp_inst_818_dout[11]),
  .I1(ram16sdp_inst_826_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1449 (
  .O(mux_o_1449),
  .I0(ram16sdp_inst_834_dout[11]),
  .I1(ram16sdp_inst_842_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1450 (
  .O(mux_o_1450),
  .I0(ram16sdp_inst_850_dout[11]),
  .I1(ram16sdp_inst_858_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1451 (
  .O(mux_o_1451),
  .I0(ram16sdp_inst_866_dout[11]),
  .I1(ram16sdp_inst_874_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1452 (
  .O(mux_o_1452),
  .I0(ram16sdp_inst_882_dout[11]),
  .I1(ram16sdp_inst_890_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1453 (
  .O(mux_o_1453),
  .I0(ram16sdp_inst_898_dout[11]),
  .I1(ram16sdp_inst_906_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1454 (
  .O(mux_o_1454),
  .I0(ram16sdp_inst_914_dout[11]),
  .I1(ram16sdp_inst_922_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1455 (
  .O(mux_o_1455),
  .I0(ram16sdp_inst_930_dout[11]),
  .I1(ram16sdp_inst_938_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1456 (
  .O(mux_o_1456),
  .I0(ram16sdp_inst_946_dout[11]),
  .I1(ram16sdp_inst_954_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1457 (
  .O(mux_o_1457),
  .I0(ram16sdp_inst_962_dout[11]),
  .I1(ram16sdp_inst_970_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1458 (
  .O(mux_o_1458),
  .I0(ram16sdp_inst_978_dout[11]),
  .I1(ram16sdp_inst_986_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1459 (
  .O(mux_o_1459),
  .I0(ram16sdp_inst_994_dout[11]),
  .I1(ram16sdp_inst_1002_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1460 (
  .O(mux_o_1460),
  .I0(ram16sdp_inst_1010_dout[11]),
  .I1(ram16sdp_inst_1018_dout[11]),
  .S0(rad[4])
);
MUX2 mux_inst_1461 (
  .O(mux_o_1461),
  .I0(mux_o_1397),
  .I1(mux_o_1398),
  .S0(rad[5])
);
MUX2 mux_inst_1462 (
  .O(mux_o_1462),
  .I0(mux_o_1399),
  .I1(mux_o_1400),
  .S0(rad[5])
);
MUX2 mux_inst_1463 (
  .O(mux_o_1463),
  .I0(mux_o_1401),
  .I1(mux_o_1402),
  .S0(rad[5])
);
MUX2 mux_inst_1464 (
  .O(mux_o_1464),
  .I0(mux_o_1403),
  .I1(mux_o_1404),
  .S0(rad[5])
);
MUX2 mux_inst_1465 (
  .O(mux_o_1465),
  .I0(mux_o_1405),
  .I1(mux_o_1406),
  .S0(rad[5])
);
MUX2 mux_inst_1466 (
  .O(mux_o_1466),
  .I0(mux_o_1407),
  .I1(mux_o_1408),
  .S0(rad[5])
);
MUX2 mux_inst_1467 (
  .O(mux_o_1467),
  .I0(mux_o_1409),
  .I1(mux_o_1410),
  .S0(rad[5])
);
MUX2 mux_inst_1468 (
  .O(mux_o_1468),
  .I0(mux_o_1411),
  .I1(mux_o_1412),
  .S0(rad[5])
);
MUX2 mux_inst_1469 (
  .O(mux_o_1469),
  .I0(mux_o_1413),
  .I1(mux_o_1414),
  .S0(rad[5])
);
MUX2 mux_inst_1470 (
  .O(mux_o_1470),
  .I0(mux_o_1415),
  .I1(mux_o_1416),
  .S0(rad[5])
);
MUX2 mux_inst_1471 (
  .O(mux_o_1471),
  .I0(mux_o_1417),
  .I1(mux_o_1418),
  .S0(rad[5])
);
MUX2 mux_inst_1472 (
  .O(mux_o_1472),
  .I0(mux_o_1419),
  .I1(mux_o_1420),
  .S0(rad[5])
);
MUX2 mux_inst_1473 (
  .O(mux_o_1473),
  .I0(mux_o_1421),
  .I1(mux_o_1422),
  .S0(rad[5])
);
MUX2 mux_inst_1474 (
  .O(mux_o_1474),
  .I0(mux_o_1423),
  .I1(mux_o_1424),
  .S0(rad[5])
);
MUX2 mux_inst_1475 (
  .O(mux_o_1475),
  .I0(mux_o_1425),
  .I1(mux_o_1426),
  .S0(rad[5])
);
MUX2 mux_inst_1476 (
  .O(mux_o_1476),
  .I0(mux_o_1427),
  .I1(mux_o_1428),
  .S0(rad[5])
);
MUX2 mux_inst_1477 (
  .O(mux_o_1477),
  .I0(mux_o_1429),
  .I1(mux_o_1430),
  .S0(rad[5])
);
MUX2 mux_inst_1478 (
  .O(mux_o_1478),
  .I0(mux_o_1431),
  .I1(mux_o_1432),
  .S0(rad[5])
);
MUX2 mux_inst_1479 (
  .O(mux_o_1479),
  .I0(mux_o_1433),
  .I1(mux_o_1434),
  .S0(rad[5])
);
MUX2 mux_inst_1480 (
  .O(mux_o_1480),
  .I0(mux_o_1435),
  .I1(mux_o_1436),
  .S0(rad[5])
);
MUX2 mux_inst_1481 (
  .O(mux_o_1481),
  .I0(mux_o_1437),
  .I1(mux_o_1438),
  .S0(rad[5])
);
MUX2 mux_inst_1482 (
  .O(mux_o_1482),
  .I0(mux_o_1439),
  .I1(mux_o_1440),
  .S0(rad[5])
);
MUX2 mux_inst_1483 (
  .O(mux_o_1483),
  .I0(mux_o_1441),
  .I1(mux_o_1442),
  .S0(rad[5])
);
MUX2 mux_inst_1484 (
  .O(mux_o_1484),
  .I0(mux_o_1443),
  .I1(mux_o_1444),
  .S0(rad[5])
);
MUX2 mux_inst_1485 (
  .O(mux_o_1485),
  .I0(mux_o_1445),
  .I1(mux_o_1446),
  .S0(rad[5])
);
MUX2 mux_inst_1486 (
  .O(mux_o_1486),
  .I0(mux_o_1447),
  .I1(mux_o_1448),
  .S0(rad[5])
);
MUX2 mux_inst_1487 (
  .O(mux_o_1487),
  .I0(mux_o_1449),
  .I1(mux_o_1450),
  .S0(rad[5])
);
MUX2 mux_inst_1488 (
  .O(mux_o_1488),
  .I0(mux_o_1451),
  .I1(mux_o_1452),
  .S0(rad[5])
);
MUX2 mux_inst_1489 (
  .O(mux_o_1489),
  .I0(mux_o_1453),
  .I1(mux_o_1454),
  .S0(rad[5])
);
MUX2 mux_inst_1490 (
  .O(mux_o_1490),
  .I0(mux_o_1455),
  .I1(mux_o_1456),
  .S0(rad[5])
);
MUX2 mux_inst_1491 (
  .O(mux_o_1491),
  .I0(mux_o_1457),
  .I1(mux_o_1458),
  .S0(rad[5])
);
MUX2 mux_inst_1492 (
  .O(mux_o_1492),
  .I0(mux_o_1459),
  .I1(mux_o_1460),
  .S0(rad[5])
);
MUX2 mux_inst_1493 (
  .O(mux_o_1493),
  .I0(mux_o_1461),
  .I1(mux_o_1462),
  .S0(rad[6])
);
MUX2 mux_inst_1494 (
  .O(mux_o_1494),
  .I0(mux_o_1463),
  .I1(mux_o_1464),
  .S0(rad[6])
);
MUX2 mux_inst_1495 (
  .O(mux_o_1495),
  .I0(mux_o_1465),
  .I1(mux_o_1466),
  .S0(rad[6])
);
MUX2 mux_inst_1496 (
  .O(mux_o_1496),
  .I0(mux_o_1467),
  .I1(mux_o_1468),
  .S0(rad[6])
);
MUX2 mux_inst_1497 (
  .O(mux_o_1497),
  .I0(mux_o_1469),
  .I1(mux_o_1470),
  .S0(rad[6])
);
MUX2 mux_inst_1498 (
  .O(mux_o_1498),
  .I0(mux_o_1471),
  .I1(mux_o_1472),
  .S0(rad[6])
);
MUX2 mux_inst_1499 (
  .O(mux_o_1499),
  .I0(mux_o_1473),
  .I1(mux_o_1474),
  .S0(rad[6])
);
MUX2 mux_inst_1500 (
  .O(mux_o_1500),
  .I0(mux_o_1475),
  .I1(mux_o_1476),
  .S0(rad[6])
);
MUX2 mux_inst_1501 (
  .O(mux_o_1501),
  .I0(mux_o_1477),
  .I1(mux_o_1478),
  .S0(rad[6])
);
MUX2 mux_inst_1502 (
  .O(mux_o_1502),
  .I0(mux_o_1479),
  .I1(mux_o_1480),
  .S0(rad[6])
);
MUX2 mux_inst_1503 (
  .O(mux_o_1503),
  .I0(mux_o_1481),
  .I1(mux_o_1482),
  .S0(rad[6])
);
MUX2 mux_inst_1504 (
  .O(mux_o_1504),
  .I0(mux_o_1483),
  .I1(mux_o_1484),
  .S0(rad[6])
);
MUX2 mux_inst_1505 (
  .O(mux_o_1505),
  .I0(mux_o_1485),
  .I1(mux_o_1486),
  .S0(rad[6])
);
MUX2 mux_inst_1506 (
  .O(mux_o_1506),
  .I0(mux_o_1487),
  .I1(mux_o_1488),
  .S0(rad[6])
);
MUX2 mux_inst_1507 (
  .O(mux_o_1507),
  .I0(mux_o_1489),
  .I1(mux_o_1490),
  .S0(rad[6])
);
MUX2 mux_inst_1508 (
  .O(mux_o_1508),
  .I0(mux_o_1491),
  .I1(mux_o_1492),
  .S0(rad[6])
);
MUX2 mux_inst_1509 (
  .O(mux_o_1509),
  .I0(mux_o_1493),
  .I1(mux_o_1494),
  .S0(rad[7])
);
MUX2 mux_inst_1510 (
  .O(mux_o_1510),
  .I0(mux_o_1495),
  .I1(mux_o_1496),
  .S0(rad[7])
);
MUX2 mux_inst_1511 (
  .O(mux_o_1511),
  .I0(mux_o_1497),
  .I1(mux_o_1498),
  .S0(rad[7])
);
MUX2 mux_inst_1512 (
  .O(mux_o_1512),
  .I0(mux_o_1499),
  .I1(mux_o_1500),
  .S0(rad[7])
);
MUX2 mux_inst_1513 (
  .O(mux_o_1513),
  .I0(mux_o_1501),
  .I1(mux_o_1502),
  .S0(rad[7])
);
MUX2 mux_inst_1514 (
  .O(mux_o_1514),
  .I0(mux_o_1503),
  .I1(mux_o_1504),
  .S0(rad[7])
);
MUX2 mux_inst_1515 (
  .O(mux_o_1515),
  .I0(mux_o_1505),
  .I1(mux_o_1506),
  .S0(rad[7])
);
MUX2 mux_inst_1516 (
  .O(mux_o_1516),
  .I0(mux_o_1507),
  .I1(mux_o_1508),
  .S0(rad[7])
);
MUX2 mux_inst_1517 (
  .O(mux_o_1517),
  .I0(mux_o_1509),
  .I1(mux_o_1510),
  .S0(rad[8])
);
MUX2 mux_inst_1518 (
  .O(mux_o_1518),
  .I0(mux_o_1511),
  .I1(mux_o_1512),
  .S0(rad[8])
);
MUX2 mux_inst_1519 (
  .O(mux_o_1519),
  .I0(mux_o_1513),
  .I1(mux_o_1514),
  .S0(rad[8])
);
MUX2 mux_inst_1520 (
  .O(mux_o_1520),
  .I0(mux_o_1515),
  .I1(mux_o_1516),
  .S0(rad[8])
);
MUX2 mux_inst_1521 (
  .O(mux_o_1521),
  .I0(mux_o_1517),
  .I1(mux_o_1518),
  .S0(rad[9])
);
MUX2 mux_inst_1522 (
  .O(mux_o_1522),
  .I0(mux_o_1519),
  .I1(mux_o_1520),
  .S0(rad[9])
);
MUX2 mux_inst_1523 (
  .O(dout[11]),
  .I0(mux_o_1521),
  .I1(mux_o_1522),
  .S0(rad[10])
);
MUX2 mux_inst_1524 (
  .O(mux_o_1524),
  .I0(ram16sdp_inst_3_dout[12]),
  .I1(ram16sdp_inst_11_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1525 (
  .O(mux_o_1525),
  .I0(ram16sdp_inst_19_dout[12]),
  .I1(ram16sdp_inst_27_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1526 (
  .O(mux_o_1526),
  .I0(ram16sdp_inst_35_dout[12]),
  .I1(ram16sdp_inst_43_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1527 (
  .O(mux_o_1527),
  .I0(ram16sdp_inst_51_dout[12]),
  .I1(ram16sdp_inst_59_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1528 (
  .O(mux_o_1528),
  .I0(ram16sdp_inst_67_dout[12]),
  .I1(ram16sdp_inst_75_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1529 (
  .O(mux_o_1529),
  .I0(ram16sdp_inst_83_dout[12]),
  .I1(ram16sdp_inst_91_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1530 (
  .O(mux_o_1530),
  .I0(ram16sdp_inst_99_dout[12]),
  .I1(ram16sdp_inst_107_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1531 (
  .O(mux_o_1531),
  .I0(ram16sdp_inst_115_dout[12]),
  .I1(ram16sdp_inst_123_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1532 (
  .O(mux_o_1532),
  .I0(ram16sdp_inst_131_dout[12]),
  .I1(ram16sdp_inst_139_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1533 (
  .O(mux_o_1533),
  .I0(ram16sdp_inst_147_dout[12]),
  .I1(ram16sdp_inst_155_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1534 (
  .O(mux_o_1534),
  .I0(ram16sdp_inst_163_dout[12]),
  .I1(ram16sdp_inst_171_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1535 (
  .O(mux_o_1535),
  .I0(ram16sdp_inst_179_dout[12]),
  .I1(ram16sdp_inst_187_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1536 (
  .O(mux_o_1536),
  .I0(ram16sdp_inst_195_dout[12]),
  .I1(ram16sdp_inst_203_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1537 (
  .O(mux_o_1537),
  .I0(ram16sdp_inst_211_dout[12]),
  .I1(ram16sdp_inst_219_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1538 (
  .O(mux_o_1538),
  .I0(ram16sdp_inst_227_dout[12]),
  .I1(ram16sdp_inst_235_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1539 (
  .O(mux_o_1539),
  .I0(ram16sdp_inst_243_dout[12]),
  .I1(ram16sdp_inst_251_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1540 (
  .O(mux_o_1540),
  .I0(ram16sdp_inst_259_dout[12]),
  .I1(ram16sdp_inst_267_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1541 (
  .O(mux_o_1541),
  .I0(ram16sdp_inst_275_dout[12]),
  .I1(ram16sdp_inst_283_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1542 (
  .O(mux_o_1542),
  .I0(ram16sdp_inst_291_dout[12]),
  .I1(ram16sdp_inst_299_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1543 (
  .O(mux_o_1543),
  .I0(ram16sdp_inst_307_dout[12]),
  .I1(ram16sdp_inst_315_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1544 (
  .O(mux_o_1544),
  .I0(ram16sdp_inst_323_dout[12]),
  .I1(ram16sdp_inst_331_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1545 (
  .O(mux_o_1545),
  .I0(ram16sdp_inst_339_dout[12]),
  .I1(ram16sdp_inst_347_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1546 (
  .O(mux_o_1546),
  .I0(ram16sdp_inst_355_dout[12]),
  .I1(ram16sdp_inst_363_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1547 (
  .O(mux_o_1547),
  .I0(ram16sdp_inst_371_dout[12]),
  .I1(ram16sdp_inst_379_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1548 (
  .O(mux_o_1548),
  .I0(ram16sdp_inst_387_dout[12]),
  .I1(ram16sdp_inst_395_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1549 (
  .O(mux_o_1549),
  .I0(ram16sdp_inst_403_dout[12]),
  .I1(ram16sdp_inst_411_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1550 (
  .O(mux_o_1550),
  .I0(ram16sdp_inst_419_dout[12]),
  .I1(ram16sdp_inst_427_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1551 (
  .O(mux_o_1551),
  .I0(ram16sdp_inst_435_dout[12]),
  .I1(ram16sdp_inst_443_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1552 (
  .O(mux_o_1552),
  .I0(ram16sdp_inst_451_dout[12]),
  .I1(ram16sdp_inst_459_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1553 (
  .O(mux_o_1553),
  .I0(ram16sdp_inst_467_dout[12]),
  .I1(ram16sdp_inst_475_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1554 (
  .O(mux_o_1554),
  .I0(ram16sdp_inst_483_dout[12]),
  .I1(ram16sdp_inst_491_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1555 (
  .O(mux_o_1555),
  .I0(ram16sdp_inst_499_dout[12]),
  .I1(ram16sdp_inst_507_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1556 (
  .O(mux_o_1556),
  .I0(ram16sdp_inst_515_dout[12]),
  .I1(ram16sdp_inst_523_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1557 (
  .O(mux_o_1557),
  .I0(ram16sdp_inst_531_dout[12]),
  .I1(ram16sdp_inst_539_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1558 (
  .O(mux_o_1558),
  .I0(ram16sdp_inst_547_dout[12]),
  .I1(ram16sdp_inst_555_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1559 (
  .O(mux_o_1559),
  .I0(ram16sdp_inst_563_dout[12]),
  .I1(ram16sdp_inst_571_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1560 (
  .O(mux_o_1560),
  .I0(ram16sdp_inst_579_dout[12]),
  .I1(ram16sdp_inst_587_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1561 (
  .O(mux_o_1561),
  .I0(ram16sdp_inst_595_dout[12]),
  .I1(ram16sdp_inst_603_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1562 (
  .O(mux_o_1562),
  .I0(ram16sdp_inst_611_dout[12]),
  .I1(ram16sdp_inst_619_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1563 (
  .O(mux_o_1563),
  .I0(ram16sdp_inst_627_dout[12]),
  .I1(ram16sdp_inst_635_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1564 (
  .O(mux_o_1564),
  .I0(ram16sdp_inst_643_dout[12]),
  .I1(ram16sdp_inst_651_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1565 (
  .O(mux_o_1565),
  .I0(ram16sdp_inst_659_dout[12]),
  .I1(ram16sdp_inst_667_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1566 (
  .O(mux_o_1566),
  .I0(ram16sdp_inst_675_dout[12]),
  .I1(ram16sdp_inst_683_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1567 (
  .O(mux_o_1567),
  .I0(ram16sdp_inst_691_dout[12]),
  .I1(ram16sdp_inst_699_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1568 (
  .O(mux_o_1568),
  .I0(ram16sdp_inst_707_dout[12]),
  .I1(ram16sdp_inst_715_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1569 (
  .O(mux_o_1569),
  .I0(ram16sdp_inst_723_dout[12]),
  .I1(ram16sdp_inst_731_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1570 (
  .O(mux_o_1570),
  .I0(ram16sdp_inst_739_dout[12]),
  .I1(ram16sdp_inst_747_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1571 (
  .O(mux_o_1571),
  .I0(ram16sdp_inst_755_dout[12]),
  .I1(ram16sdp_inst_763_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1572 (
  .O(mux_o_1572),
  .I0(ram16sdp_inst_771_dout[12]),
  .I1(ram16sdp_inst_779_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1573 (
  .O(mux_o_1573),
  .I0(ram16sdp_inst_787_dout[12]),
  .I1(ram16sdp_inst_795_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1574 (
  .O(mux_o_1574),
  .I0(ram16sdp_inst_803_dout[12]),
  .I1(ram16sdp_inst_811_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1575 (
  .O(mux_o_1575),
  .I0(ram16sdp_inst_819_dout[12]),
  .I1(ram16sdp_inst_827_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1576 (
  .O(mux_o_1576),
  .I0(ram16sdp_inst_835_dout[12]),
  .I1(ram16sdp_inst_843_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1577 (
  .O(mux_o_1577),
  .I0(ram16sdp_inst_851_dout[12]),
  .I1(ram16sdp_inst_859_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1578 (
  .O(mux_o_1578),
  .I0(ram16sdp_inst_867_dout[12]),
  .I1(ram16sdp_inst_875_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1579 (
  .O(mux_o_1579),
  .I0(ram16sdp_inst_883_dout[12]),
  .I1(ram16sdp_inst_891_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1580 (
  .O(mux_o_1580),
  .I0(ram16sdp_inst_899_dout[12]),
  .I1(ram16sdp_inst_907_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1581 (
  .O(mux_o_1581),
  .I0(ram16sdp_inst_915_dout[12]),
  .I1(ram16sdp_inst_923_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1582 (
  .O(mux_o_1582),
  .I0(ram16sdp_inst_931_dout[12]),
  .I1(ram16sdp_inst_939_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1583 (
  .O(mux_o_1583),
  .I0(ram16sdp_inst_947_dout[12]),
  .I1(ram16sdp_inst_955_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1584 (
  .O(mux_o_1584),
  .I0(ram16sdp_inst_963_dout[12]),
  .I1(ram16sdp_inst_971_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1585 (
  .O(mux_o_1585),
  .I0(ram16sdp_inst_979_dout[12]),
  .I1(ram16sdp_inst_987_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1586 (
  .O(mux_o_1586),
  .I0(ram16sdp_inst_995_dout[12]),
  .I1(ram16sdp_inst_1003_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1587 (
  .O(mux_o_1587),
  .I0(ram16sdp_inst_1011_dout[12]),
  .I1(ram16sdp_inst_1019_dout[12]),
  .S0(rad[4])
);
MUX2 mux_inst_1588 (
  .O(mux_o_1588),
  .I0(mux_o_1524),
  .I1(mux_o_1525),
  .S0(rad[5])
);
MUX2 mux_inst_1589 (
  .O(mux_o_1589),
  .I0(mux_o_1526),
  .I1(mux_o_1527),
  .S0(rad[5])
);
MUX2 mux_inst_1590 (
  .O(mux_o_1590),
  .I0(mux_o_1528),
  .I1(mux_o_1529),
  .S0(rad[5])
);
MUX2 mux_inst_1591 (
  .O(mux_o_1591),
  .I0(mux_o_1530),
  .I1(mux_o_1531),
  .S0(rad[5])
);
MUX2 mux_inst_1592 (
  .O(mux_o_1592),
  .I0(mux_o_1532),
  .I1(mux_o_1533),
  .S0(rad[5])
);
MUX2 mux_inst_1593 (
  .O(mux_o_1593),
  .I0(mux_o_1534),
  .I1(mux_o_1535),
  .S0(rad[5])
);
MUX2 mux_inst_1594 (
  .O(mux_o_1594),
  .I0(mux_o_1536),
  .I1(mux_o_1537),
  .S0(rad[5])
);
MUX2 mux_inst_1595 (
  .O(mux_o_1595),
  .I0(mux_o_1538),
  .I1(mux_o_1539),
  .S0(rad[5])
);
MUX2 mux_inst_1596 (
  .O(mux_o_1596),
  .I0(mux_o_1540),
  .I1(mux_o_1541),
  .S0(rad[5])
);
MUX2 mux_inst_1597 (
  .O(mux_o_1597),
  .I0(mux_o_1542),
  .I1(mux_o_1543),
  .S0(rad[5])
);
MUX2 mux_inst_1598 (
  .O(mux_o_1598),
  .I0(mux_o_1544),
  .I1(mux_o_1545),
  .S0(rad[5])
);
MUX2 mux_inst_1599 (
  .O(mux_o_1599),
  .I0(mux_o_1546),
  .I1(mux_o_1547),
  .S0(rad[5])
);
MUX2 mux_inst_1600 (
  .O(mux_o_1600),
  .I0(mux_o_1548),
  .I1(mux_o_1549),
  .S0(rad[5])
);
MUX2 mux_inst_1601 (
  .O(mux_o_1601),
  .I0(mux_o_1550),
  .I1(mux_o_1551),
  .S0(rad[5])
);
MUX2 mux_inst_1602 (
  .O(mux_o_1602),
  .I0(mux_o_1552),
  .I1(mux_o_1553),
  .S0(rad[5])
);
MUX2 mux_inst_1603 (
  .O(mux_o_1603),
  .I0(mux_o_1554),
  .I1(mux_o_1555),
  .S0(rad[5])
);
MUX2 mux_inst_1604 (
  .O(mux_o_1604),
  .I0(mux_o_1556),
  .I1(mux_o_1557),
  .S0(rad[5])
);
MUX2 mux_inst_1605 (
  .O(mux_o_1605),
  .I0(mux_o_1558),
  .I1(mux_o_1559),
  .S0(rad[5])
);
MUX2 mux_inst_1606 (
  .O(mux_o_1606),
  .I0(mux_o_1560),
  .I1(mux_o_1561),
  .S0(rad[5])
);
MUX2 mux_inst_1607 (
  .O(mux_o_1607),
  .I0(mux_o_1562),
  .I1(mux_o_1563),
  .S0(rad[5])
);
MUX2 mux_inst_1608 (
  .O(mux_o_1608),
  .I0(mux_o_1564),
  .I1(mux_o_1565),
  .S0(rad[5])
);
MUX2 mux_inst_1609 (
  .O(mux_o_1609),
  .I0(mux_o_1566),
  .I1(mux_o_1567),
  .S0(rad[5])
);
MUX2 mux_inst_1610 (
  .O(mux_o_1610),
  .I0(mux_o_1568),
  .I1(mux_o_1569),
  .S0(rad[5])
);
MUX2 mux_inst_1611 (
  .O(mux_o_1611),
  .I0(mux_o_1570),
  .I1(mux_o_1571),
  .S0(rad[5])
);
MUX2 mux_inst_1612 (
  .O(mux_o_1612),
  .I0(mux_o_1572),
  .I1(mux_o_1573),
  .S0(rad[5])
);
MUX2 mux_inst_1613 (
  .O(mux_o_1613),
  .I0(mux_o_1574),
  .I1(mux_o_1575),
  .S0(rad[5])
);
MUX2 mux_inst_1614 (
  .O(mux_o_1614),
  .I0(mux_o_1576),
  .I1(mux_o_1577),
  .S0(rad[5])
);
MUX2 mux_inst_1615 (
  .O(mux_o_1615),
  .I0(mux_o_1578),
  .I1(mux_o_1579),
  .S0(rad[5])
);
MUX2 mux_inst_1616 (
  .O(mux_o_1616),
  .I0(mux_o_1580),
  .I1(mux_o_1581),
  .S0(rad[5])
);
MUX2 mux_inst_1617 (
  .O(mux_o_1617),
  .I0(mux_o_1582),
  .I1(mux_o_1583),
  .S0(rad[5])
);
MUX2 mux_inst_1618 (
  .O(mux_o_1618),
  .I0(mux_o_1584),
  .I1(mux_o_1585),
  .S0(rad[5])
);
MUX2 mux_inst_1619 (
  .O(mux_o_1619),
  .I0(mux_o_1586),
  .I1(mux_o_1587),
  .S0(rad[5])
);
MUX2 mux_inst_1620 (
  .O(mux_o_1620),
  .I0(mux_o_1588),
  .I1(mux_o_1589),
  .S0(rad[6])
);
MUX2 mux_inst_1621 (
  .O(mux_o_1621),
  .I0(mux_o_1590),
  .I1(mux_o_1591),
  .S0(rad[6])
);
MUX2 mux_inst_1622 (
  .O(mux_o_1622),
  .I0(mux_o_1592),
  .I1(mux_o_1593),
  .S0(rad[6])
);
MUX2 mux_inst_1623 (
  .O(mux_o_1623),
  .I0(mux_o_1594),
  .I1(mux_o_1595),
  .S0(rad[6])
);
MUX2 mux_inst_1624 (
  .O(mux_o_1624),
  .I0(mux_o_1596),
  .I1(mux_o_1597),
  .S0(rad[6])
);
MUX2 mux_inst_1625 (
  .O(mux_o_1625),
  .I0(mux_o_1598),
  .I1(mux_o_1599),
  .S0(rad[6])
);
MUX2 mux_inst_1626 (
  .O(mux_o_1626),
  .I0(mux_o_1600),
  .I1(mux_o_1601),
  .S0(rad[6])
);
MUX2 mux_inst_1627 (
  .O(mux_o_1627),
  .I0(mux_o_1602),
  .I1(mux_o_1603),
  .S0(rad[6])
);
MUX2 mux_inst_1628 (
  .O(mux_o_1628),
  .I0(mux_o_1604),
  .I1(mux_o_1605),
  .S0(rad[6])
);
MUX2 mux_inst_1629 (
  .O(mux_o_1629),
  .I0(mux_o_1606),
  .I1(mux_o_1607),
  .S0(rad[6])
);
MUX2 mux_inst_1630 (
  .O(mux_o_1630),
  .I0(mux_o_1608),
  .I1(mux_o_1609),
  .S0(rad[6])
);
MUX2 mux_inst_1631 (
  .O(mux_o_1631),
  .I0(mux_o_1610),
  .I1(mux_o_1611),
  .S0(rad[6])
);
MUX2 mux_inst_1632 (
  .O(mux_o_1632),
  .I0(mux_o_1612),
  .I1(mux_o_1613),
  .S0(rad[6])
);
MUX2 mux_inst_1633 (
  .O(mux_o_1633),
  .I0(mux_o_1614),
  .I1(mux_o_1615),
  .S0(rad[6])
);
MUX2 mux_inst_1634 (
  .O(mux_o_1634),
  .I0(mux_o_1616),
  .I1(mux_o_1617),
  .S0(rad[6])
);
MUX2 mux_inst_1635 (
  .O(mux_o_1635),
  .I0(mux_o_1618),
  .I1(mux_o_1619),
  .S0(rad[6])
);
MUX2 mux_inst_1636 (
  .O(mux_o_1636),
  .I0(mux_o_1620),
  .I1(mux_o_1621),
  .S0(rad[7])
);
MUX2 mux_inst_1637 (
  .O(mux_o_1637),
  .I0(mux_o_1622),
  .I1(mux_o_1623),
  .S0(rad[7])
);
MUX2 mux_inst_1638 (
  .O(mux_o_1638),
  .I0(mux_o_1624),
  .I1(mux_o_1625),
  .S0(rad[7])
);
MUX2 mux_inst_1639 (
  .O(mux_o_1639),
  .I0(mux_o_1626),
  .I1(mux_o_1627),
  .S0(rad[7])
);
MUX2 mux_inst_1640 (
  .O(mux_o_1640),
  .I0(mux_o_1628),
  .I1(mux_o_1629),
  .S0(rad[7])
);
MUX2 mux_inst_1641 (
  .O(mux_o_1641),
  .I0(mux_o_1630),
  .I1(mux_o_1631),
  .S0(rad[7])
);
MUX2 mux_inst_1642 (
  .O(mux_o_1642),
  .I0(mux_o_1632),
  .I1(mux_o_1633),
  .S0(rad[7])
);
MUX2 mux_inst_1643 (
  .O(mux_o_1643),
  .I0(mux_o_1634),
  .I1(mux_o_1635),
  .S0(rad[7])
);
MUX2 mux_inst_1644 (
  .O(mux_o_1644),
  .I0(mux_o_1636),
  .I1(mux_o_1637),
  .S0(rad[8])
);
MUX2 mux_inst_1645 (
  .O(mux_o_1645),
  .I0(mux_o_1638),
  .I1(mux_o_1639),
  .S0(rad[8])
);
MUX2 mux_inst_1646 (
  .O(mux_o_1646),
  .I0(mux_o_1640),
  .I1(mux_o_1641),
  .S0(rad[8])
);
MUX2 mux_inst_1647 (
  .O(mux_o_1647),
  .I0(mux_o_1642),
  .I1(mux_o_1643),
  .S0(rad[8])
);
MUX2 mux_inst_1648 (
  .O(mux_o_1648),
  .I0(mux_o_1644),
  .I1(mux_o_1645),
  .S0(rad[9])
);
MUX2 mux_inst_1649 (
  .O(mux_o_1649),
  .I0(mux_o_1646),
  .I1(mux_o_1647),
  .S0(rad[9])
);
MUX2 mux_inst_1650 (
  .O(dout[12]),
  .I0(mux_o_1648),
  .I1(mux_o_1649),
  .S0(rad[10])
);
MUX2 mux_inst_1651 (
  .O(mux_o_1651),
  .I0(ram16sdp_inst_3_dout[13]),
  .I1(ram16sdp_inst_11_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1652 (
  .O(mux_o_1652),
  .I0(ram16sdp_inst_19_dout[13]),
  .I1(ram16sdp_inst_27_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1653 (
  .O(mux_o_1653),
  .I0(ram16sdp_inst_35_dout[13]),
  .I1(ram16sdp_inst_43_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1654 (
  .O(mux_o_1654),
  .I0(ram16sdp_inst_51_dout[13]),
  .I1(ram16sdp_inst_59_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1655 (
  .O(mux_o_1655),
  .I0(ram16sdp_inst_67_dout[13]),
  .I1(ram16sdp_inst_75_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1656 (
  .O(mux_o_1656),
  .I0(ram16sdp_inst_83_dout[13]),
  .I1(ram16sdp_inst_91_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1657 (
  .O(mux_o_1657),
  .I0(ram16sdp_inst_99_dout[13]),
  .I1(ram16sdp_inst_107_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1658 (
  .O(mux_o_1658),
  .I0(ram16sdp_inst_115_dout[13]),
  .I1(ram16sdp_inst_123_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1659 (
  .O(mux_o_1659),
  .I0(ram16sdp_inst_131_dout[13]),
  .I1(ram16sdp_inst_139_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1660 (
  .O(mux_o_1660),
  .I0(ram16sdp_inst_147_dout[13]),
  .I1(ram16sdp_inst_155_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1661 (
  .O(mux_o_1661),
  .I0(ram16sdp_inst_163_dout[13]),
  .I1(ram16sdp_inst_171_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1662 (
  .O(mux_o_1662),
  .I0(ram16sdp_inst_179_dout[13]),
  .I1(ram16sdp_inst_187_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1663 (
  .O(mux_o_1663),
  .I0(ram16sdp_inst_195_dout[13]),
  .I1(ram16sdp_inst_203_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1664 (
  .O(mux_o_1664),
  .I0(ram16sdp_inst_211_dout[13]),
  .I1(ram16sdp_inst_219_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1665 (
  .O(mux_o_1665),
  .I0(ram16sdp_inst_227_dout[13]),
  .I1(ram16sdp_inst_235_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1666 (
  .O(mux_o_1666),
  .I0(ram16sdp_inst_243_dout[13]),
  .I1(ram16sdp_inst_251_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1667 (
  .O(mux_o_1667),
  .I0(ram16sdp_inst_259_dout[13]),
  .I1(ram16sdp_inst_267_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1668 (
  .O(mux_o_1668),
  .I0(ram16sdp_inst_275_dout[13]),
  .I1(ram16sdp_inst_283_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1669 (
  .O(mux_o_1669),
  .I0(ram16sdp_inst_291_dout[13]),
  .I1(ram16sdp_inst_299_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1670 (
  .O(mux_o_1670),
  .I0(ram16sdp_inst_307_dout[13]),
  .I1(ram16sdp_inst_315_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1671 (
  .O(mux_o_1671),
  .I0(ram16sdp_inst_323_dout[13]),
  .I1(ram16sdp_inst_331_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1672 (
  .O(mux_o_1672),
  .I0(ram16sdp_inst_339_dout[13]),
  .I1(ram16sdp_inst_347_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1673 (
  .O(mux_o_1673),
  .I0(ram16sdp_inst_355_dout[13]),
  .I1(ram16sdp_inst_363_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1674 (
  .O(mux_o_1674),
  .I0(ram16sdp_inst_371_dout[13]),
  .I1(ram16sdp_inst_379_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1675 (
  .O(mux_o_1675),
  .I0(ram16sdp_inst_387_dout[13]),
  .I1(ram16sdp_inst_395_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1676 (
  .O(mux_o_1676),
  .I0(ram16sdp_inst_403_dout[13]),
  .I1(ram16sdp_inst_411_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1677 (
  .O(mux_o_1677),
  .I0(ram16sdp_inst_419_dout[13]),
  .I1(ram16sdp_inst_427_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1678 (
  .O(mux_o_1678),
  .I0(ram16sdp_inst_435_dout[13]),
  .I1(ram16sdp_inst_443_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1679 (
  .O(mux_o_1679),
  .I0(ram16sdp_inst_451_dout[13]),
  .I1(ram16sdp_inst_459_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1680 (
  .O(mux_o_1680),
  .I0(ram16sdp_inst_467_dout[13]),
  .I1(ram16sdp_inst_475_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1681 (
  .O(mux_o_1681),
  .I0(ram16sdp_inst_483_dout[13]),
  .I1(ram16sdp_inst_491_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1682 (
  .O(mux_o_1682),
  .I0(ram16sdp_inst_499_dout[13]),
  .I1(ram16sdp_inst_507_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1683 (
  .O(mux_o_1683),
  .I0(ram16sdp_inst_515_dout[13]),
  .I1(ram16sdp_inst_523_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1684 (
  .O(mux_o_1684),
  .I0(ram16sdp_inst_531_dout[13]),
  .I1(ram16sdp_inst_539_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1685 (
  .O(mux_o_1685),
  .I0(ram16sdp_inst_547_dout[13]),
  .I1(ram16sdp_inst_555_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1686 (
  .O(mux_o_1686),
  .I0(ram16sdp_inst_563_dout[13]),
  .I1(ram16sdp_inst_571_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1687 (
  .O(mux_o_1687),
  .I0(ram16sdp_inst_579_dout[13]),
  .I1(ram16sdp_inst_587_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1688 (
  .O(mux_o_1688),
  .I0(ram16sdp_inst_595_dout[13]),
  .I1(ram16sdp_inst_603_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1689 (
  .O(mux_o_1689),
  .I0(ram16sdp_inst_611_dout[13]),
  .I1(ram16sdp_inst_619_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1690 (
  .O(mux_o_1690),
  .I0(ram16sdp_inst_627_dout[13]),
  .I1(ram16sdp_inst_635_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1691 (
  .O(mux_o_1691),
  .I0(ram16sdp_inst_643_dout[13]),
  .I1(ram16sdp_inst_651_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1692 (
  .O(mux_o_1692),
  .I0(ram16sdp_inst_659_dout[13]),
  .I1(ram16sdp_inst_667_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1693 (
  .O(mux_o_1693),
  .I0(ram16sdp_inst_675_dout[13]),
  .I1(ram16sdp_inst_683_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1694 (
  .O(mux_o_1694),
  .I0(ram16sdp_inst_691_dout[13]),
  .I1(ram16sdp_inst_699_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1695 (
  .O(mux_o_1695),
  .I0(ram16sdp_inst_707_dout[13]),
  .I1(ram16sdp_inst_715_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1696 (
  .O(mux_o_1696),
  .I0(ram16sdp_inst_723_dout[13]),
  .I1(ram16sdp_inst_731_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1697 (
  .O(mux_o_1697),
  .I0(ram16sdp_inst_739_dout[13]),
  .I1(ram16sdp_inst_747_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1698 (
  .O(mux_o_1698),
  .I0(ram16sdp_inst_755_dout[13]),
  .I1(ram16sdp_inst_763_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1699 (
  .O(mux_o_1699),
  .I0(ram16sdp_inst_771_dout[13]),
  .I1(ram16sdp_inst_779_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1700 (
  .O(mux_o_1700),
  .I0(ram16sdp_inst_787_dout[13]),
  .I1(ram16sdp_inst_795_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1701 (
  .O(mux_o_1701),
  .I0(ram16sdp_inst_803_dout[13]),
  .I1(ram16sdp_inst_811_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1702 (
  .O(mux_o_1702),
  .I0(ram16sdp_inst_819_dout[13]),
  .I1(ram16sdp_inst_827_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1703 (
  .O(mux_o_1703),
  .I0(ram16sdp_inst_835_dout[13]),
  .I1(ram16sdp_inst_843_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1704 (
  .O(mux_o_1704),
  .I0(ram16sdp_inst_851_dout[13]),
  .I1(ram16sdp_inst_859_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1705 (
  .O(mux_o_1705),
  .I0(ram16sdp_inst_867_dout[13]),
  .I1(ram16sdp_inst_875_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1706 (
  .O(mux_o_1706),
  .I0(ram16sdp_inst_883_dout[13]),
  .I1(ram16sdp_inst_891_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1707 (
  .O(mux_o_1707),
  .I0(ram16sdp_inst_899_dout[13]),
  .I1(ram16sdp_inst_907_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1708 (
  .O(mux_o_1708),
  .I0(ram16sdp_inst_915_dout[13]),
  .I1(ram16sdp_inst_923_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1709 (
  .O(mux_o_1709),
  .I0(ram16sdp_inst_931_dout[13]),
  .I1(ram16sdp_inst_939_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1710 (
  .O(mux_o_1710),
  .I0(ram16sdp_inst_947_dout[13]),
  .I1(ram16sdp_inst_955_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1711 (
  .O(mux_o_1711),
  .I0(ram16sdp_inst_963_dout[13]),
  .I1(ram16sdp_inst_971_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1712 (
  .O(mux_o_1712),
  .I0(ram16sdp_inst_979_dout[13]),
  .I1(ram16sdp_inst_987_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1713 (
  .O(mux_o_1713),
  .I0(ram16sdp_inst_995_dout[13]),
  .I1(ram16sdp_inst_1003_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1714 (
  .O(mux_o_1714),
  .I0(ram16sdp_inst_1011_dout[13]),
  .I1(ram16sdp_inst_1019_dout[13]),
  .S0(rad[4])
);
MUX2 mux_inst_1715 (
  .O(mux_o_1715),
  .I0(mux_o_1651),
  .I1(mux_o_1652),
  .S0(rad[5])
);
MUX2 mux_inst_1716 (
  .O(mux_o_1716),
  .I0(mux_o_1653),
  .I1(mux_o_1654),
  .S0(rad[5])
);
MUX2 mux_inst_1717 (
  .O(mux_o_1717),
  .I0(mux_o_1655),
  .I1(mux_o_1656),
  .S0(rad[5])
);
MUX2 mux_inst_1718 (
  .O(mux_o_1718),
  .I0(mux_o_1657),
  .I1(mux_o_1658),
  .S0(rad[5])
);
MUX2 mux_inst_1719 (
  .O(mux_o_1719),
  .I0(mux_o_1659),
  .I1(mux_o_1660),
  .S0(rad[5])
);
MUX2 mux_inst_1720 (
  .O(mux_o_1720),
  .I0(mux_o_1661),
  .I1(mux_o_1662),
  .S0(rad[5])
);
MUX2 mux_inst_1721 (
  .O(mux_o_1721),
  .I0(mux_o_1663),
  .I1(mux_o_1664),
  .S0(rad[5])
);
MUX2 mux_inst_1722 (
  .O(mux_o_1722),
  .I0(mux_o_1665),
  .I1(mux_o_1666),
  .S0(rad[5])
);
MUX2 mux_inst_1723 (
  .O(mux_o_1723),
  .I0(mux_o_1667),
  .I1(mux_o_1668),
  .S0(rad[5])
);
MUX2 mux_inst_1724 (
  .O(mux_o_1724),
  .I0(mux_o_1669),
  .I1(mux_o_1670),
  .S0(rad[5])
);
MUX2 mux_inst_1725 (
  .O(mux_o_1725),
  .I0(mux_o_1671),
  .I1(mux_o_1672),
  .S0(rad[5])
);
MUX2 mux_inst_1726 (
  .O(mux_o_1726),
  .I0(mux_o_1673),
  .I1(mux_o_1674),
  .S0(rad[5])
);
MUX2 mux_inst_1727 (
  .O(mux_o_1727),
  .I0(mux_o_1675),
  .I1(mux_o_1676),
  .S0(rad[5])
);
MUX2 mux_inst_1728 (
  .O(mux_o_1728),
  .I0(mux_o_1677),
  .I1(mux_o_1678),
  .S0(rad[5])
);
MUX2 mux_inst_1729 (
  .O(mux_o_1729),
  .I0(mux_o_1679),
  .I1(mux_o_1680),
  .S0(rad[5])
);
MUX2 mux_inst_1730 (
  .O(mux_o_1730),
  .I0(mux_o_1681),
  .I1(mux_o_1682),
  .S0(rad[5])
);
MUX2 mux_inst_1731 (
  .O(mux_o_1731),
  .I0(mux_o_1683),
  .I1(mux_o_1684),
  .S0(rad[5])
);
MUX2 mux_inst_1732 (
  .O(mux_o_1732),
  .I0(mux_o_1685),
  .I1(mux_o_1686),
  .S0(rad[5])
);
MUX2 mux_inst_1733 (
  .O(mux_o_1733),
  .I0(mux_o_1687),
  .I1(mux_o_1688),
  .S0(rad[5])
);
MUX2 mux_inst_1734 (
  .O(mux_o_1734),
  .I0(mux_o_1689),
  .I1(mux_o_1690),
  .S0(rad[5])
);
MUX2 mux_inst_1735 (
  .O(mux_o_1735),
  .I0(mux_o_1691),
  .I1(mux_o_1692),
  .S0(rad[5])
);
MUX2 mux_inst_1736 (
  .O(mux_o_1736),
  .I0(mux_o_1693),
  .I1(mux_o_1694),
  .S0(rad[5])
);
MUX2 mux_inst_1737 (
  .O(mux_o_1737),
  .I0(mux_o_1695),
  .I1(mux_o_1696),
  .S0(rad[5])
);
MUX2 mux_inst_1738 (
  .O(mux_o_1738),
  .I0(mux_o_1697),
  .I1(mux_o_1698),
  .S0(rad[5])
);
MUX2 mux_inst_1739 (
  .O(mux_o_1739),
  .I0(mux_o_1699),
  .I1(mux_o_1700),
  .S0(rad[5])
);
MUX2 mux_inst_1740 (
  .O(mux_o_1740),
  .I0(mux_o_1701),
  .I1(mux_o_1702),
  .S0(rad[5])
);
MUX2 mux_inst_1741 (
  .O(mux_o_1741),
  .I0(mux_o_1703),
  .I1(mux_o_1704),
  .S0(rad[5])
);
MUX2 mux_inst_1742 (
  .O(mux_o_1742),
  .I0(mux_o_1705),
  .I1(mux_o_1706),
  .S0(rad[5])
);
MUX2 mux_inst_1743 (
  .O(mux_o_1743),
  .I0(mux_o_1707),
  .I1(mux_o_1708),
  .S0(rad[5])
);
MUX2 mux_inst_1744 (
  .O(mux_o_1744),
  .I0(mux_o_1709),
  .I1(mux_o_1710),
  .S0(rad[5])
);
MUX2 mux_inst_1745 (
  .O(mux_o_1745),
  .I0(mux_o_1711),
  .I1(mux_o_1712),
  .S0(rad[5])
);
MUX2 mux_inst_1746 (
  .O(mux_o_1746),
  .I0(mux_o_1713),
  .I1(mux_o_1714),
  .S0(rad[5])
);
MUX2 mux_inst_1747 (
  .O(mux_o_1747),
  .I0(mux_o_1715),
  .I1(mux_o_1716),
  .S0(rad[6])
);
MUX2 mux_inst_1748 (
  .O(mux_o_1748),
  .I0(mux_o_1717),
  .I1(mux_o_1718),
  .S0(rad[6])
);
MUX2 mux_inst_1749 (
  .O(mux_o_1749),
  .I0(mux_o_1719),
  .I1(mux_o_1720),
  .S0(rad[6])
);
MUX2 mux_inst_1750 (
  .O(mux_o_1750),
  .I0(mux_o_1721),
  .I1(mux_o_1722),
  .S0(rad[6])
);
MUX2 mux_inst_1751 (
  .O(mux_o_1751),
  .I0(mux_o_1723),
  .I1(mux_o_1724),
  .S0(rad[6])
);
MUX2 mux_inst_1752 (
  .O(mux_o_1752),
  .I0(mux_o_1725),
  .I1(mux_o_1726),
  .S0(rad[6])
);
MUX2 mux_inst_1753 (
  .O(mux_o_1753),
  .I0(mux_o_1727),
  .I1(mux_o_1728),
  .S0(rad[6])
);
MUX2 mux_inst_1754 (
  .O(mux_o_1754),
  .I0(mux_o_1729),
  .I1(mux_o_1730),
  .S0(rad[6])
);
MUX2 mux_inst_1755 (
  .O(mux_o_1755),
  .I0(mux_o_1731),
  .I1(mux_o_1732),
  .S0(rad[6])
);
MUX2 mux_inst_1756 (
  .O(mux_o_1756),
  .I0(mux_o_1733),
  .I1(mux_o_1734),
  .S0(rad[6])
);
MUX2 mux_inst_1757 (
  .O(mux_o_1757),
  .I0(mux_o_1735),
  .I1(mux_o_1736),
  .S0(rad[6])
);
MUX2 mux_inst_1758 (
  .O(mux_o_1758),
  .I0(mux_o_1737),
  .I1(mux_o_1738),
  .S0(rad[6])
);
MUX2 mux_inst_1759 (
  .O(mux_o_1759),
  .I0(mux_o_1739),
  .I1(mux_o_1740),
  .S0(rad[6])
);
MUX2 mux_inst_1760 (
  .O(mux_o_1760),
  .I0(mux_o_1741),
  .I1(mux_o_1742),
  .S0(rad[6])
);
MUX2 mux_inst_1761 (
  .O(mux_o_1761),
  .I0(mux_o_1743),
  .I1(mux_o_1744),
  .S0(rad[6])
);
MUX2 mux_inst_1762 (
  .O(mux_o_1762),
  .I0(mux_o_1745),
  .I1(mux_o_1746),
  .S0(rad[6])
);
MUX2 mux_inst_1763 (
  .O(mux_o_1763),
  .I0(mux_o_1747),
  .I1(mux_o_1748),
  .S0(rad[7])
);
MUX2 mux_inst_1764 (
  .O(mux_o_1764),
  .I0(mux_o_1749),
  .I1(mux_o_1750),
  .S0(rad[7])
);
MUX2 mux_inst_1765 (
  .O(mux_o_1765),
  .I0(mux_o_1751),
  .I1(mux_o_1752),
  .S0(rad[7])
);
MUX2 mux_inst_1766 (
  .O(mux_o_1766),
  .I0(mux_o_1753),
  .I1(mux_o_1754),
  .S0(rad[7])
);
MUX2 mux_inst_1767 (
  .O(mux_o_1767),
  .I0(mux_o_1755),
  .I1(mux_o_1756),
  .S0(rad[7])
);
MUX2 mux_inst_1768 (
  .O(mux_o_1768),
  .I0(mux_o_1757),
  .I1(mux_o_1758),
  .S0(rad[7])
);
MUX2 mux_inst_1769 (
  .O(mux_o_1769),
  .I0(mux_o_1759),
  .I1(mux_o_1760),
  .S0(rad[7])
);
MUX2 mux_inst_1770 (
  .O(mux_o_1770),
  .I0(mux_o_1761),
  .I1(mux_o_1762),
  .S0(rad[7])
);
MUX2 mux_inst_1771 (
  .O(mux_o_1771),
  .I0(mux_o_1763),
  .I1(mux_o_1764),
  .S0(rad[8])
);
MUX2 mux_inst_1772 (
  .O(mux_o_1772),
  .I0(mux_o_1765),
  .I1(mux_o_1766),
  .S0(rad[8])
);
MUX2 mux_inst_1773 (
  .O(mux_o_1773),
  .I0(mux_o_1767),
  .I1(mux_o_1768),
  .S0(rad[8])
);
MUX2 mux_inst_1774 (
  .O(mux_o_1774),
  .I0(mux_o_1769),
  .I1(mux_o_1770),
  .S0(rad[8])
);
MUX2 mux_inst_1775 (
  .O(mux_o_1775),
  .I0(mux_o_1771),
  .I1(mux_o_1772),
  .S0(rad[9])
);
MUX2 mux_inst_1776 (
  .O(mux_o_1776),
  .I0(mux_o_1773),
  .I1(mux_o_1774),
  .S0(rad[9])
);
MUX2 mux_inst_1777 (
  .O(dout[13]),
  .I0(mux_o_1775),
  .I1(mux_o_1776),
  .S0(rad[10])
);
MUX2 mux_inst_1778 (
  .O(mux_o_1778),
  .I0(ram16sdp_inst_3_dout[14]),
  .I1(ram16sdp_inst_11_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1779 (
  .O(mux_o_1779),
  .I0(ram16sdp_inst_19_dout[14]),
  .I1(ram16sdp_inst_27_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1780 (
  .O(mux_o_1780),
  .I0(ram16sdp_inst_35_dout[14]),
  .I1(ram16sdp_inst_43_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1781 (
  .O(mux_o_1781),
  .I0(ram16sdp_inst_51_dout[14]),
  .I1(ram16sdp_inst_59_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1782 (
  .O(mux_o_1782),
  .I0(ram16sdp_inst_67_dout[14]),
  .I1(ram16sdp_inst_75_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1783 (
  .O(mux_o_1783),
  .I0(ram16sdp_inst_83_dout[14]),
  .I1(ram16sdp_inst_91_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1784 (
  .O(mux_o_1784),
  .I0(ram16sdp_inst_99_dout[14]),
  .I1(ram16sdp_inst_107_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1785 (
  .O(mux_o_1785),
  .I0(ram16sdp_inst_115_dout[14]),
  .I1(ram16sdp_inst_123_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1786 (
  .O(mux_o_1786),
  .I0(ram16sdp_inst_131_dout[14]),
  .I1(ram16sdp_inst_139_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1787 (
  .O(mux_o_1787),
  .I0(ram16sdp_inst_147_dout[14]),
  .I1(ram16sdp_inst_155_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1788 (
  .O(mux_o_1788),
  .I0(ram16sdp_inst_163_dout[14]),
  .I1(ram16sdp_inst_171_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1789 (
  .O(mux_o_1789),
  .I0(ram16sdp_inst_179_dout[14]),
  .I1(ram16sdp_inst_187_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1790 (
  .O(mux_o_1790),
  .I0(ram16sdp_inst_195_dout[14]),
  .I1(ram16sdp_inst_203_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1791 (
  .O(mux_o_1791),
  .I0(ram16sdp_inst_211_dout[14]),
  .I1(ram16sdp_inst_219_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1792 (
  .O(mux_o_1792),
  .I0(ram16sdp_inst_227_dout[14]),
  .I1(ram16sdp_inst_235_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1793 (
  .O(mux_o_1793),
  .I0(ram16sdp_inst_243_dout[14]),
  .I1(ram16sdp_inst_251_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1794 (
  .O(mux_o_1794),
  .I0(ram16sdp_inst_259_dout[14]),
  .I1(ram16sdp_inst_267_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1795 (
  .O(mux_o_1795),
  .I0(ram16sdp_inst_275_dout[14]),
  .I1(ram16sdp_inst_283_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1796 (
  .O(mux_o_1796),
  .I0(ram16sdp_inst_291_dout[14]),
  .I1(ram16sdp_inst_299_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1797 (
  .O(mux_o_1797),
  .I0(ram16sdp_inst_307_dout[14]),
  .I1(ram16sdp_inst_315_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1798 (
  .O(mux_o_1798),
  .I0(ram16sdp_inst_323_dout[14]),
  .I1(ram16sdp_inst_331_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1799 (
  .O(mux_o_1799),
  .I0(ram16sdp_inst_339_dout[14]),
  .I1(ram16sdp_inst_347_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1800 (
  .O(mux_o_1800),
  .I0(ram16sdp_inst_355_dout[14]),
  .I1(ram16sdp_inst_363_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1801 (
  .O(mux_o_1801),
  .I0(ram16sdp_inst_371_dout[14]),
  .I1(ram16sdp_inst_379_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1802 (
  .O(mux_o_1802),
  .I0(ram16sdp_inst_387_dout[14]),
  .I1(ram16sdp_inst_395_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1803 (
  .O(mux_o_1803),
  .I0(ram16sdp_inst_403_dout[14]),
  .I1(ram16sdp_inst_411_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1804 (
  .O(mux_o_1804),
  .I0(ram16sdp_inst_419_dout[14]),
  .I1(ram16sdp_inst_427_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1805 (
  .O(mux_o_1805),
  .I0(ram16sdp_inst_435_dout[14]),
  .I1(ram16sdp_inst_443_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1806 (
  .O(mux_o_1806),
  .I0(ram16sdp_inst_451_dout[14]),
  .I1(ram16sdp_inst_459_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1807 (
  .O(mux_o_1807),
  .I0(ram16sdp_inst_467_dout[14]),
  .I1(ram16sdp_inst_475_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1808 (
  .O(mux_o_1808),
  .I0(ram16sdp_inst_483_dout[14]),
  .I1(ram16sdp_inst_491_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1809 (
  .O(mux_o_1809),
  .I0(ram16sdp_inst_499_dout[14]),
  .I1(ram16sdp_inst_507_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1810 (
  .O(mux_o_1810),
  .I0(ram16sdp_inst_515_dout[14]),
  .I1(ram16sdp_inst_523_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1811 (
  .O(mux_o_1811),
  .I0(ram16sdp_inst_531_dout[14]),
  .I1(ram16sdp_inst_539_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1812 (
  .O(mux_o_1812),
  .I0(ram16sdp_inst_547_dout[14]),
  .I1(ram16sdp_inst_555_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1813 (
  .O(mux_o_1813),
  .I0(ram16sdp_inst_563_dout[14]),
  .I1(ram16sdp_inst_571_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1814 (
  .O(mux_o_1814),
  .I0(ram16sdp_inst_579_dout[14]),
  .I1(ram16sdp_inst_587_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1815 (
  .O(mux_o_1815),
  .I0(ram16sdp_inst_595_dout[14]),
  .I1(ram16sdp_inst_603_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1816 (
  .O(mux_o_1816),
  .I0(ram16sdp_inst_611_dout[14]),
  .I1(ram16sdp_inst_619_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1817 (
  .O(mux_o_1817),
  .I0(ram16sdp_inst_627_dout[14]),
  .I1(ram16sdp_inst_635_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1818 (
  .O(mux_o_1818),
  .I0(ram16sdp_inst_643_dout[14]),
  .I1(ram16sdp_inst_651_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1819 (
  .O(mux_o_1819),
  .I0(ram16sdp_inst_659_dout[14]),
  .I1(ram16sdp_inst_667_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1820 (
  .O(mux_o_1820),
  .I0(ram16sdp_inst_675_dout[14]),
  .I1(ram16sdp_inst_683_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1821 (
  .O(mux_o_1821),
  .I0(ram16sdp_inst_691_dout[14]),
  .I1(ram16sdp_inst_699_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1822 (
  .O(mux_o_1822),
  .I0(ram16sdp_inst_707_dout[14]),
  .I1(ram16sdp_inst_715_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1823 (
  .O(mux_o_1823),
  .I0(ram16sdp_inst_723_dout[14]),
  .I1(ram16sdp_inst_731_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1824 (
  .O(mux_o_1824),
  .I0(ram16sdp_inst_739_dout[14]),
  .I1(ram16sdp_inst_747_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1825 (
  .O(mux_o_1825),
  .I0(ram16sdp_inst_755_dout[14]),
  .I1(ram16sdp_inst_763_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1826 (
  .O(mux_o_1826),
  .I0(ram16sdp_inst_771_dout[14]),
  .I1(ram16sdp_inst_779_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1827 (
  .O(mux_o_1827),
  .I0(ram16sdp_inst_787_dout[14]),
  .I1(ram16sdp_inst_795_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1828 (
  .O(mux_o_1828),
  .I0(ram16sdp_inst_803_dout[14]),
  .I1(ram16sdp_inst_811_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1829 (
  .O(mux_o_1829),
  .I0(ram16sdp_inst_819_dout[14]),
  .I1(ram16sdp_inst_827_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1830 (
  .O(mux_o_1830),
  .I0(ram16sdp_inst_835_dout[14]),
  .I1(ram16sdp_inst_843_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1831 (
  .O(mux_o_1831),
  .I0(ram16sdp_inst_851_dout[14]),
  .I1(ram16sdp_inst_859_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1832 (
  .O(mux_o_1832),
  .I0(ram16sdp_inst_867_dout[14]),
  .I1(ram16sdp_inst_875_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1833 (
  .O(mux_o_1833),
  .I0(ram16sdp_inst_883_dout[14]),
  .I1(ram16sdp_inst_891_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1834 (
  .O(mux_o_1834),
  .I0(ram16sdp_inst_899_dout[14]),
  .I1(ram16sdp_inst_907_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1835 (
  .O(mux_o_1835),
  .I0(ram16sdp_inst_915_dout[14]),
  .I1(ram16sdp_inst_923_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1836 (
  .O(mux_o_1836),
  .I0(ram16sdp_inst_931_dout[14]),
  .I1(ram16sdp_inst_939_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1837 (
  .O(mux_o_1837),
  .I0(ram16sdp_inst_947_dout[14]),
  .I1(ram16sdp_inst_955_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1838 (
  .O(mux_o_1838),
  .I0(ram16sdp_inst_963_dout[14]),
  .I1(ram16sdp_inst_971_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1839 (
  .O(mux_o_1839),
  .I0(ram16sdp_inst_979_dout[14]),
  .I1(ram16sdp_inst_987_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1840 (
  .O(mux_o_1840),
  .I0(ram16sdp_inst_995_dout[14]),
  .I1(ram16sdp_inst_1003_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1841 (
  .O(mux_o_1841),
  .I0(ram16sdp_inst_1011_dout[14]),
  .I1(ram16sdp_inst_1019_dout[14]),
  .S0(rad[4])
);
MUX2 mux_inst_1842 (
  .O(mux_o_1842),
  .I0(mux_o_1778),
  .I1(mux_o_1779),
  .S0(rad[5])
);
MUX2 mux_inst_1843 (
  .O(mux_o_1843),
  .I0(mux_o_1780),
  .I1(mux_o_1781),
  .S0(rad[5])
);
MUX2 mux_inst_1844 (
  .O(mux_o_1844),
  .I0(mux_o_1782),
  .I1(mux_o_1783),
  .S0(rad[5])
);
MUX2 mux_inst_1845 (
  .O(mux_o_1845),
  .I0(mux_o_1784),
  .I1(mux_o_1785),
  .S0(rad[5])
);
MUX2 mux_inst_1846 (
  .O(mux_o_1846),
  .I0(mux_o_1786),
  .I1(mux_o_1787),
  .S0(rad[5])
);
MUX2 mux_inst_1847 (
  .O(mux_o_1847),
  .I0(mux_o_1788),
  .I1(mux_o_1789),
  .S0(rad[5])
);
MUX2 mux_inst_1848 (
  .O(mux_o_1848),
  .I0(mux_o_1790),
  .I1(mux_o_1791),
  .S0(rad[5])
);
MUX2 mux_inst_1849 (
  .O(mux_o_1849),
  .I0(mux_o_1792),
  .I1(mux_o_1793),
  .S0(rad[5])
);
MUX2 mux_inst_1850 (
  .O(mux_o_1850),
  .I0(mux_o_1794),
  .I1(mux_o_1795),
  .S0(rad[5])
);
MUX2 mux_inst_1851 (
  .O(mux_o_1851),
  .I0(mux_o_1796),
  .I1(mux_o_1797),
  .S0(rad[5])
);
MUX2 mux_inst_1852 (
  .O(mux_o_1852),
  .I0(mux_o_1798),
  .I1(mux_o_1799),
  .S0(rad[5])
);
MUX2 mux_inst_1853 (
  .O(mux_o_1853),
  .I0(mux_o_1800),
  .I1(mux_o_1801),
  .S0(rad[5])
);
MUX2 mux_inst_1854 (
  .O(mux_o_1854),
  .I0(mux_o_1802),
  .I1(mux_o_1803),
  .S0(rad[5])
);
MUX2 mux_inst_1855 (
  .O(mux_o_1855),
  .I0(mux_o_1804),
  .I1(mux_o_1805),
  .S0(rad[5])
);
MUX2 mux_inst_1856 (
  .O(mux_o_1856),
  .I0(mux_o_1806),
  .I1(mux_o_1807),
  .S0(rad[5])
);
MUX2 mux_inst_1857 (
  .O(mux_o_1857),
  .I0(mux_o_1808),
  .I1(mux_o_1809),
  .S0(rad[5])
);
MUX2 mux_inst_1858 (
  .O(mux_o_1858),
  .I0(mux_o_1810),
  .I1(mux_o_1811),
  .S0(rad[5])
);
MUX2 mux_inst_1859 (
  .O(mux_o_1859),
  .I0(mux_o_1812),
  .I1(mux_o_1813),
  .S0(rad[5])
);
MUX2 mux_inst_1860 (
  .O(mux_o_1860),
  .I0(mux_o_1814),
  .I1(mux_o_1815),
  .S0(rad[5])
);
MUX2 mux_inst_1861 (
  .O(mux_o_1861),
  .I0(mux_o_1816),
  .I1(mux_o_1817),
  .S0(rad[5])
);
MUX2 mux_inst_1862 (
  .O(mux_o_1862),
  .I0(mux_o_1818),
  .I1(mux_o_1819),
  .S0(rad[5])
);
MUX2 mux_inst_1863 (
  .O(mux_o_1863),
  .I0(mux_o_1820),
  .I1(mux_o_1821),
  .S0(rad[5])
);
MUX2 mux_inst_1864 (
  .O(mux_o_1864),
  .I0(mux_o_1822),
  .I1(mux_o_1823),
  .S0(rad[5])
);
MUX2 mux_inst_1865 (
  .O(mux_o_1865),
  .I0(mux_o_1824),
  .I1(mux_o_1825),
  .S0(rad[5])
);
MUX2 mux_inst_1866 (
  .O(mux_o_1866),
  .I0(mux_o_1826),
  .I1(mux_o_1827),
  .S0(rad[5])
);
MUX2 mux_inst_1867 (
  .O(mux_o_1867),
  .I0(mux_o_1828),
  .I1(mux_o_1829),
  .S0(rad[5])
);
MUX2 mux_inst_1868 (
  .O(mux_o_1868),
  .I0(mux_o_1830),
  .I1(mux_o_1831),
  .S0(rad[5])
);
MUX2 mux_inst_1869 (
  .O(mux_o_1869),
  .I0(mux_o_1832),
  .I1(mux_o_1833),
  .S0(rad[5])
);
MUX2 mux_inst_1870 (
  .O(mux_o_1870),
  .I0(mux_o_1834),
  .I1(mux_o_1835),
  .S0(rad[5])
);
MUX2 mux_inst_1871 (
  .O(mux_o_1871),
  .I0(mux_o_1836),
  .I1(mux_o_1837),
  .S0(rad[5])
);
MUX2 mux_inst_1872 (
  .O(mux_o_1872),
  .I0(mux_o_1838),
  .I1(mux_o_1839),
  .S0(rad[5])
);
MUX2 mux_inst_1873 (
  .O(mux_o_1873),
  .I0(mux_o_1840),
  .I1(mux_o_1841),
  .S0(rad[5])
);
MUX2 mux_inst_1874 (
  .O(mux_o_1874),
  .I0(mux_o_1842),
  .I1(mux_o_1843),
  .S0(rad[6])
);
MUX2 mux_inst_1875 (
  .O(mux_o_1875),
  .I0(mux_o_1844),
  .I1(mux_o_1845),
  .S0(rad[6])
);
MUX2 mux_inst_1876 (
  .O(mux_o_1876),
  .I0(mux_o_1846),
  .I1(mux_o_1847),
  .S0(rad[6])
);
MUX2 mux_inst_1877 (
  .O(mux_o_1877),
  .I0(mux_o_1848),
  .I1(mux_o_1849),
  .S0(rad[6])
);
MUX2 mux_inst_1878 (
  .O(mux_o_1878),
  .I0(mux_o_1850),
  .I1(mux_o_1851),
  .S0(rad[6])
);
MUX2 mux_inst_1879 (
  .O(mux_o_1879),
  .I0(mux_o_1852),
  .I1(mux_o_1853),
  .S0(rad[6])
);
MUX2 mux_inst_1880 (
  .O(mux_o_1880),
  .I0(mux_o_1854),
  .I1(mux_o_1855),
  .S0(rad[6])
);
MUX2 mux_inst_1881 (
  .O(mux_o_1881),
  .I0(mux_o_1856),
  .I1(mux_o_1857),
  .S0(rad[6])
);
MUX2 mux_inst_1882 (
  .O(mux_o_1882),
  .I0(mux_o_1858),
  .I1(mux_o_1859),
  .S0(rad[6])
);
MUX2 mux_inst_1883 (
  .O(mux_o_1883),
  .I0(mux_o_1860),
  .I1(mux_o_1861),
  .S0(rad[6])
);
MUX2 mux_inst_1884 (
  .O(mux_o_1884),
  .I0(mux_o_1862),
  .I1(mux_o_1863),
  .S0(rad[6])
);
MUX2 mux_inst_1885 (
  .O(mux_o_1885),
  .I0(mux_o_1864),
  .I1(mux_o_1865),
  .S0(rad[6])
);
MUX2 mux_inst_1886 (
  .O(mux_o_1886),
  .I0(mux_o_1866),
  .I1(mux_o_1867),
  .S0(rad[6])
);
MUX2 mux_inst_1887 (
  .O(mux_o_1887),
  .I0(mux_o_1868),
  .I1(mux_o_1869),
  .S0(rad[6])
);
MUX2 mux_inst_1888 (
  .O(mux_o_1888),
  .I0(mux_o_1870),
  .I1(mux_o_1871),
  .S0(rad[6])
);
MUX2 mux_inst_1889 (
  .O(mux_o_1889),
  .I0(mux_o_1872),
  .I1(mux_o_1873),
  .S0(rad[6])
);
MUX2 mux_inst_1890 (
  .O(mux_o_1890),
  .I0(mux_o_1874),
  .I1(mux_o_1875),
  .S0(rad[7])
);
MUX2 mux_inst_1891 (
  .O(mux_o_1891),
  .I0(mux_o_1876),
  .I1(mux_o_1877),
  .S0(rad[7])
);
MUX2 mux_inst_1892 (
  .O(mux_o_1892),
  .I0(mux_o_1878),
  .I1(mux_o_1879),
  .S0(rad[7])
);
MUX2 mux_inst_1893 (
  .O(mux_o_1893),
  .I0(mux_o_1880),
  .I1(mux_o_1881),
  .S0(rad[7])
);
MUX2 mux_inst_1894 (
  .O(mux_o_1894),
  .I0(mux_o_1882),
  .I1(mux_o_1883),
  .S0(rad[7])
);
MUX2 mux_inst_1895 (
  .O(mux_o_1895),
  .I0(mux_o_1884),
  .I1(mux_o_1885),
  .S0(rad[7])
);
MUX2 mux_inst_1896 (
  .O(mux_o_1896),
  .I0(mux_o_1886),
  .I1(mux_o_1887),
  .S0(rad[7])
);
MUX2 mux_inst_1897 (
  .O(mux_o_1897),
  .I0(mux_o_1888),
  .I1(mux_o_1889),
  .S0(rad[7])
);
MUX2 mux_inst_1898 (
  .O(mux_o_1898),
  .I0(mux_o_1890),
  .I1(mux_o_1891),
  .S0(rad[8])
);
MUX2 mux_inst_1899 (
  .O(mux_o_1899),
  .I0(mux_o_1892),
  .I1(mux_o_1893),
  .S0(rad[8])
);
MUX2 mux_inst_1900 (
  .O(mux_o_1900),
  .I0(mux_o_1894),
  .I1(mux_o_1895),
  .S0(rad[8])
);
MUX2 mux_inst_1901 (
  .O(mux_o_1901),
  .I0(mux_o_1896),
  .I1(mux_o_1897),
  .S0(rad[8])
);
MUX2 mux_inst_1902 (
  .O(mux_o_1902),
  .I0(mux_o_1898),
  .I1(mux_o_1899),
  .S0(rad[9])
);
MUX2 mux_inst_1903 (
  .O(mux_o_1903),
  .I0(mux_o_1900),
  .I1(mux_o_1901),
  .S0(rad[9])
);
MUX2 mux_inst_1904 (
  .O(dout[14]),
  .I0(mux_o_1902),
  .I1(mux_o_1903),
  .S0(rad[10])
);
MUX2 mux_inst_1905 (
  .O(mux_o_1905),
  .I0(ram16sdp_inst_3_dout[15]),
  .I1(ram16sdp_inst_11_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1906 (
  .O(mux_o_1906),
  .I0(ram16sdp_inst_19_dout[15]),
  .I1(ram16sdp_inst_27_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1907 (
  .O(mux_o_1907),
  .I0(ram16sdp_inst_35_dout[15]),
  .I1(ram16sdp_inst_43_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1908 (
  .O(mux_o_1908),
  .I0(ram16sdp_inst_51_dout[15]),
  .I1(ram16sdp_inst_59_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1909 (
  .O(mux_o_1909),
  .I0(ram16sdp_inst_67_dout[15]),
  .I1(ram16sdp_inst_75_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1910 (
  .O(mux_o_1910),
  .I0(ram16sdp_inst_83_dout[15]),
  .I1(ram16sdp_inst_91_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1911 (
  .O(mux_o_1911),
  .I0(ram16sdp_inst_99_dout[15]),
  .I1(ram16sdp_inst_107_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1912 (
  .O(mux_o_1912),
  .I0(ram16sdp_inst_115_dout[15]),
  .I1(ram16sdp_inst_123_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1913 (
  .O(mux_o_1913),
  .I0(ram16sdp_inst_131_dout[15]),
  .I1(ram16sdp_inst_139_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1914 (
  .O(mux_o_1914),
  .I0(ram16sdp_inst_147_dout[15]),
  .I1(ram16sdp_inst_155_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1915 (
  .O(mux_o_1915),
  .I0(ram16sdp_inst_163_dout[15]),
  .I1(ram16sdp_inst_171_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1916 (
  .O(mux_o_1916),
  .I0(ram16sdp_inst_179_dout[15]),
  .I1(ram16sdp_inst_187_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1917 (
  .O(mux_o_1917),
  .I0(ram16sdp_inst_195_dout[15]),
  .I1(ram16sdp_inst_203_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1918 (
  .O(mux_o_1918),
  .I0(ram16sdp_inst_211_dout[15]),
  .I1(ram16sdp_inst_219_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1919 (
  .O(mux_o_1919),
  .I0(ram16sdp_inst_227_dout[15]),
  .I1(ram16sdp_inst_235_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1920 (
  .O(mux_o_1920),
  .I0(ram16sdp_inst_243_dout[15]),
  .I1(ram16sdp_inst_251_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1921 (
  .O(mux_o_1921),
  .I0(ram16sdp_inst_259_dout[15]),
  .I1(ram16sdp_inst_267_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1922 (
  .O(mux_o_1922),
  .I0(ram16sdp_inst_275_dout[15]),
  .I1(ram16sdp_inst_283_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1923 (
  .O(mux_o_1923),
  .I0(ram16sdp_inst_291_dout[15]),
  .I1(ram16sdp_inst_299_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1924 (
  .O(mux_o_1924),
  .I0(ram16sdp_inst_307_dout[15]),
  .I1(ram16sdp_inst_315_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1925 (
  .O(mux_o_1925),
  .I0(ram16sdp_inst_323_dout[15]),
  .I1(ram16sdp_inst_331_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1926 (
  .O(mux_o_1926),
  .I0(ram16sdp_inst_339_dout[15]),
  .I1(ram16sdp_inst_347_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1927 (
  .O(mux_o_1927),
  .I0(ram16sdp_inst_355_dout[15]),
  .I1(ram16sdp_inst_363_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1928 (
  .O(mux_o_1928),
  .I0(ram16sdp_inst_371_dout[15]),
  .I1(ram16sdp_inst_379_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1929 (
  .O(mux_o_1929),
  .I0(ram16sdp_inst_387_dout[15]),
  .I1(ram16sdp_inst_395_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1930 (
  .O(mux_o_1930),
  .I0(ram16sdp_inst_403_dout[15]),
  .I1(ram16sdp_inst_411_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1931 (
  .O(mux_o_1931),
  .I0(ram16sdp_inst_419_dout[15]),
  .I1(ram16sdp_inst_427_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1932 (
  .O(mux_o_1932),
  .I0(ram16sdp_inst_435_dout[15]),
  .I1(ram16sdp_inst_443_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1933 (
  .O(mux_o_1933),
  .I0(ram16sdp_inst_451_dout[15]),
  .I1(ram16sdp_inst_459_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1934 (
  .O(mux_o_1934),
  .I0(ram16sdp_inst_467_dout[15]),
  .I1(ram16sdp_inst_475_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1935 (
  .O(mux_o_1935),
  .I0(ram16sdp_inst_483_dout[15]),
  .I1(ram16sdp_inst_491_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1936 (
  .O(mux_o_1936),
  .I0(ram16sdp_inst_499_dout[15]),
  .I1(ram16sdp_inst_507_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1937 (
  .O(mux_o_1937),
  .I0(ram16sdp_inst_515_dout[15]),
  .I1(ram16sdp_inst_523_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1938 (
  .O(mux_o_1938),
  .I0(ram16sdp_inst_531_dout[15]),
  .I1(ram16sdp_inst_539_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1939 (
  .O(mux_o_1939),
  .I0(ram16sdp_inst_547_dout[15]),
  .I1(ram16sdp_inst_555_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1940 (
  .O(mux_o_1940),
  .I0(ram16sdp_inst_563_dout[15]),
  .I1(ram16sdp_inst_571_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1941 (
  .O(mux_o_1941),
  .I0(ram16sdp_inst_579_dout[15]),
  .I1(ram16sdp_inst_587_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1942 (
  .O(mux_o_1942),
  .I0(ram16sdp_inst_595_dout[15]),
  .I1(ram16sdp_inst_603_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1943 (
  .O(mux_o_1943),
  .I0(ram16sdp_inst_611_dout[15]),
  .I1(ram16sdp_inst_619_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1944 (
  .O(mux_o_1944),
  .I0(ram16sdp_inst_627_dout[15]),
  .I1(ram16sdp_inst_635_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1945 (
  .O(mux_o_1945),
  .I0(ram16sdp_inst_643_dout[15]),
  .I1(ram16sdp_inst_651_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1946 (
  .O(mux_o_1946),
  .I0(ram16sdp_inst_659_dout[15]),
  .I1(ram16sdp_inst_667_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1947 (
  .O(mux_o_1947),
  .I0(ram16sdp_inst_675_dout[15]),
  .I1(ram16sdp_inst_683_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1948 (
  .O(mux_o_1948),
  .I0(ram16sdp_inst_691_dout[15]),
  .I1(ram16sdp_inst_699_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1949 (
  .O(mux_o_1949),
  .I0(ram16sdp_inst_707_dout[15]),
  .I1(ram16sdp_inst_715_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1950 (
  .O(mux_o_1950),
  .I0(ram16sdp_inst_723_dout[15]),
  .I1(ram16sdp_inst_731_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1951 (
  .O(mux_o_1951),
  .I0(ram16sdp_inst_739_dout[15]),
  .I1(ram16sdp_inst_747_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1952 (
  .O(mux_o_1952),
  .I0(ram16sdp_inst_755_dout[15]),
  .I1(ram16sdp_inst_763_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1953 (
  .O(mux_o_1953),
  .I0(ram16sdp_inst_771_dout[15]),
  .I1(ram16sdp_inst_779_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1954 (
  .O(mux_o_1954),
  .I0(ram16sdp_inst_787_dout[15]),
  .I1(ram16sdp_inst_795_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1955 (
  .O(mux_o_1955),
  .I0(ram16sdp_inst_803_dout[15]),
  .I1(ram16sdp_inst_811_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1956 (
  .O(mux_o_1956),
  .I0(ram16sdp_inst_819_dout[15]),
  .I1(ram16sdp_inst_827_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1957 (
  .O(mux_o_1957),
  .I0(ram16sdp_inst_835_dout[15]),
  .I1(ram16sdp_inst_843_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1958 (
  .O(mux_o_1958),
  .I0(ram16sdp_inst_851_dout[15]),
  .I1(ram16sdp_inst_859_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1959 (
  .O(mux_o_1959),
  .I0(ram16sdp_inst_867_dout[15]),
  .I1(ram16sdp_inst_875_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1960 (
  .O(mux_o_1960),
  .I0(ram16sdp_inst_883_dout[15]),
  .I1(ram16sdp_inst_891_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1961 (
  .O(mux_o_1961),
  .I0(ram16sdp_inst_899_dout[15]),
  .I1(ram16sdp_inst_907_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1962 (
  .O(mux_o_1962),
  .I0(ram16sdp_inst_915_dout[15]),
  .I1(ram16sdp_inst_923_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1963 (
  .O(mux_o_1963),
  .I0(ram16sdp_inst_931_dout[15]),
  .I1(ram16sdp_inst_939_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1964 (
  .O(mux_o_1964),
  .I0(ram16sdp_inst_947_dout[15]),
  .I1(ram16sdp_inst_955_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1965 (
  .O(mux_o_1965),
  .I0(ram16sdp_inst_963_dout[15]),
  .I1(ram16sdp_inst_971_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1966 (
  .O(mux_o_1966),
  .I0(ram16sdp_inst_979_dout[15]),
  .I1(ram16sdp_inst_987_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1967 (
  .O(mux_o_1967),
  .I0(ram16sdp_inst_995_dout[15]),
  .I1(ram16sdp_inst_1003_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1968 (
  .O(mux_o_1968),
  .I0(ram16sdp_inst_1011_dout[15]),
  .I1(ram16sdp_inst_1019_dout[15]),
  .S0(rad[4])
);
MUX2 mux_inst_1969 (
  .O(mux_o_1969),
  .I0(mux_o_1905),
  .I1(mux_o_1906),
  .S0(rad[5])
);
MUX2 mux_inst_1970 (
  .O(mux_o_1970),
  .I0(mux_o_1907),
  .I1(mux_o_1908),
  .S0(rad[5])
);
MUX2 mux_inst_1971 (
  .O(mux_o_1971),
  .I0(mux_o_1909),
  .I1(mux_o_1910),
  .S0(rad[5])
);
MUX2 mux_inst_1972 (
  .O(mux_o_1972),
  .I0(mux_o_1911),
  .I1(mux_o_1912),
  .S0(rad[5])
);
MUX2 mux_inst_1973 (
  .O(mux_o_1973),
  .I0(mux_o_1913),
  .I1(mux_o_1914),
  .S0(rad[5])
);
MUX2 mux_inst_1974 (
  .O(mux_o_1974),
  .I0(mux_o_1915),
  .I1(mux_o_1916),
  .S0(rad[5])
);
MUX2 mux_inst_1975 (
  .O(mux_o_1975),
  .I0(mux_o_1917),
  .I1(mux_o_1918),
  .S0(rad[5])
);
MUX2 mux_inst_1976 (
  .O(mux_o_1976),
  .I0(mux_o_1919),
  .I1(mux_o_1920),
  .S0(rad[5])
);
MUX2 mux_inst_1977 (
  .O(mux_o_1977),
  .I0(mux_o_1921),
  .I1(mux_o_1922),
  .S0(rad[5])
);
MUX2 mux_inst_1978 (
  .O(mux_o_1978),
  .I0(mux_o_1923),
  .I1(mux_o_1924),
  .S0(rad[5])
);
MUX2 mux_inst_1979 (
  .O(mux_o_1979),
  .I0(mux_o_1925),
  .I1(mux_o_1926),
  .S0(rad[5])
);
MUX2 mux_inst_1980 (
  .O(mux_o_1980),
  .I0(mux_o_1927),
  .I1(mux_o_1928),
  .S0(rad[5])
);
MUX2 mux_inst_1981 (
  .O(mux_o_1981),
  .I0(mux_o_1929),
  .I1(mux_o_1930),
  .S0(rad[5])
);
MUX2 mux_inst_1982 (
  .O(mux_o_1982),
  .I0(mux_o_1931),
  .I1(mux_o_1932),
  .S0(rad[5])
);
MUX2 mux_inst_1983 (
  .O(mux_o_1983),
  .I0(mux_o_1933),
  .I1(mux_o_1934),
  .S0(rad[5])
);
MUX2 mux_inst_1984 (
  .O(mux_o_1984),
  .I0(mux_o_1935),
  .I1(mux_o_1936),
  .S0(rad[5])
);
MUX2 mux_inst_1985 (
  .O(mux_o_1985),
  .I0(mux_o_1937),
  .I1(mux_o_1938),
  .S0(rad[5])
);
MUX2 mux_inst_1986 (
  .O(mux_o_1986),
  .I0(mux_o_1939),
  .I1(mux_o_1940),
  .S0(rad[5])
);
MUX2 mux_inst_1987 (
  .O(mux_o_1987),
  .I0(mux_o_1941),
  .I1(mux_o_1942),
  .S0(rad[5])
);
MUX2 mux_inst_1988 (
  .O(mux_o_1988),
  .I0(mux_o_1943),
  .I1(mux_o_1944),
  .S0(rad[5])
);
MUX2 mux_inst_1989 (
  .O(mux_o_1989),
  .I0(mux_o_1945),
  .I1(mux_o_1946),
  .S0(rad[5])
);
MUX2 mux_inst_1990 (
  .O(mux_o_1990),
  .I0(mux_o_1947),
  .I1(mux_o_1948),
  .S0(rad[5])
);
MUX2 mux_inst_1991 (
  .O(mux_o_1991),
  .I0(mux_o_1949),
  .I1(mux_o_1950),
  .S0(rad[5])
);
MUX2 mux_inst_1992 (
  .O(mux_o_1992),
  .I0(mux_o_1951),
  .I1(mux_o_1952),
  .S0(rad[5])
);
MUX2 mux_inst_1993 (
  .O(mux_o_1993),
  .I0(mux_o_1953),
  .I1(mux_o_1954),
  .S0(rad[5])
);
MUX2 mux_inst_1994 (
  .O(mux_o_1994),
  .I0(mux_o_1955),
  .I1(mux_o_1956),
  .S0(rad[5])
);
MUX2 mux_inst_1995 (
  .O(mux_o_1995),
  .I0(mux_o_1957),
  .I1(mux_o_1958),
  .S0(rad[5])
);
MUX2 mux_inst_1996 (
  .O(mux_o_1996),
  .I0(mux_o_1959),
  .I1(mux_o_1960),
  .S0(rad[5])
);
MUX2 mux_inst_1997 (
  .O(mux_o_1997),
  .I0(mux_o_1961),
  .I1(mux_o_1962),
  .S0(rad[5])
);
MUX2 mux_inst_1998 (
  .O(mux_o_1998),
  .I0(mux_o_1963),
  .I1(mux_o_1964),
  .S0(rad[5])
);
MUX2 mux_inst_1999 (
  .O(mux_o_1999),
  .I0(mux_o_1965),
  .I1(mux_o_1966),
  .S0(rad[5])
);
MUX2 mux_inst_2000 (
  .O(mux_o_2000),
  .I0(mux_o_1967),
  .I1(mux_o_1968),
  .S0(rad[5])
);
MUX2 mux_inst_2001 (
  .O(mux_o_2001),
  .I0(mux_o_1969),
  .I1(mux_o_1970),
  .S0(rad[6])
);
MUX2 mux_inst_2002 (
  .O(mux_o_2002),
  .I0(mux_o_1971),
  .I1(mux_o_1972),
  .S0(rad[6])
);
MUX2 mux_inst_2003 (
  .O(mux_o_2003),
  .I0(mux_o_1973),
  .I1(mux_o_1974),
  .S0(rad[6])
);
MUX2 mux_inst_2004 (
  .O(mux_o_2004),
  .I0(mux_o_1975),
  .I1(mux_o_1976),
  .S0(rad[6])
);
MUX2 mux_inst_2005 (
  .O(mux_o_2005),
  .I0(mux_o_1977),
  .I1(mux_o_1978),
  .S0(rad[6])
);
MUX2 mux_inst_2006 (
  .O(mux_o_2006),
  .I0(mux_o_1979),
  .I1(mux_o_1980),
  .S0(rad[6])
);
MUX2 mux_inst_2007 (
  .O(mux_o_2007),
  .I0(mux_o_1981),
  .I1(mux_o_1982),
  .S0(rad[6])
);
MUX2 mux_inst_2008 (
  .O(mux_o_2008),
  .I0(mux_o_1983),
  .I1(mux_o_1984),
  .S0(rad[6])
);
MUX2 mux_inst_2009 (
  .O(mux_o_2009),
  .I0(mux_o_1985),
  .I1(mux_o_1986),
  .S0(rad[6])
);
MUX2 mux_inst_2010 (
  .O(mux_o_2010),
  .I0(mux_o_1987),
  .I1(mux_o_1988),
  .S0(rad[6])
);
MUX2 mux_inst_2011 (
  .O(mux_o_2011),
  .I0(mux_o_1989),
  .I1(mux_o_1990),
  .S0(rad[6])
);
MUX2 mux_inst_2012 (
  .O(mux_o_2012),
  .I0(mux_o_1991),
  .I1(mux_o_1992),
  .S0(rad[6])
);
MUX2 mux_inst_2013 (
  .O(mux_o_2013),
  .I0(mux_o_1993),
  .I1(mux_o_1994),
  .S0(rad[6])
);
MUX2 mux_inst_2014 (
  .O(mux_o_2014),
  .I0(mux_o_1995),
  .I1(mux_o_1996),
  .S0(rad[6])
);
MUX2 mux_inst_2015 (
  .O(mux_o_2015),
  .I0(mux_o_1997),
  .I1(mux_o_1998),
  .S0(rad[6])
);
MUX2 mux_inst_2016 (
  .O(mux_o_2016),
  .I0(mux_o_1999),
  .I1(mux_o_2000),
  .S0(rad[6])
);
MUX2 mux_inst_2017 (
  .O(mux_o_2017),
  .I0(mux_o_2001),
  .I1(mux_o_2002),
  .S0(rad[7])
);
MUX2 mux_inst_2018 (
  .O(mux_o_2018),
  .I0(mux_o_2003),
  .I1(mux_o_2004),
  .S0(rad[7])
);
MUX2 mux_inst_2019 (
  .O(mux_o_2019),
  .I0(mux_o_2005),
  .I1(mux_o_2006),
  .S0(rad[7])
);
MUX2 mux_inst_2020 (
  .O(mux_o_2020),
  .I0(mux_o_2007),
  .I1(mux_o_2008),
  .S0(rad[7])
);
MUX2 mux_inst_2021 (
  .O(mux_o_2021),
  .I0(mux_o_2009),
  .I1(mux_o_2010),
  .S0(rad[7])
);
MUX2 mux_inst_2022 (
  .O(mux_o_2022),
  .I0(mux_o_2011),
  .I1(mux_o_2012),
  .S0(rad[7])
);
MUX2 mux_inst_2023 (
  .O(mux_o_2023),
  .I0(mux_o_2013),
  .I1(mux_o_2014),
  .S0(rad[7])
);
MUX2 mux_inst_2024 (
  .O(mux_o_2024),
  .I0(mux_o_2015),
  .I1(mux_o_2016),
  .S0(rad[7])
);
MUX2 mux_inst_2025 (
  .O(mux_o_2025),
  .I0(mux_o_2017),
  .I1(mux_o_2018),
  .S0(rad[8])
);
MUX2 mux_inst_2026 (
  .O(mux_o_2026),
  .I0(mux_o_2019),
  .I1(mux_o_2020),
  .S0(rad[8])
);
MUX2 mux_inst_2027 (
  .O(mux_o_2027),
  .I0(mux_o_2021),
  .I1(mux_o_2022),
  .S0(rad[8])
);
MUX2 mux_inst_2028 (
  .O(mux_o_2028),
  .I0(mux_o_2023),
  .I1(mux_o_2024),
  .S0(rad[8])
);
MUX2 mux_inst_2029 (
  .O(mux_o_2029),
  .I0(mux_o_2025),
  .I1(mux_o_2026),
  .S0(rad[9])
);
MUX2 mux_inst_2030 (
  .O(mux_o_2030),
  .I0(mux_o_2027),
  .I1(mux_o_2028),
  .S0(rad[9])
);
MUX2 mux_inst_2031 (
  .O(dout[15]),
  .I0(mux_o_2029),
  .I1(mux_o_2030),
  .S0(rad[10])
);
MUX2 mux_inst_2032 (
  .O(mux_o_2032),
  .I0(ram16sdp_inst_4_dout[16]),
  .I1(ram16sdp_inst_12_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2033 (
  .O(mux_o_2033),
  .I0(ram16sdp_inst_20_dout[16]),
  .I1(ram16sdp_inst_28_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2034 (
  .O(mux_o_2034),
  .I0(ram16sdp_inst_36_dout[16]),
  .I1(ram16sdp_inst_44_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2035 (
  .O(mux_o_2035),
  .I0(ram16sdp_inst_52_dout[16]),
  .I1(ram16sdp_inst_60_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2036 (
  .O(mux_o_2036),
  .I0(ram16sdp_inst_68_dout[16]),
  .I1(ram16sdp_inst_76_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2037 (
  .O(mux_o_2037),
  .I0(ram16sdp_inst_84_dout[16]),
  .I1(ram16sdp_inst_92_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2038 (
  .O(mux_o_2038),
  .I0(ram16sdp_inst_100_dout[16]),
  .I1(ram16sdp_inst_108_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2039 (
  .O(mux_o_2039),
  .I0(ram16sdp_inst_116_dout[16]),
  .I1(ram16sdp_inst_124_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2040 (
  .O(mux_o_2040),
  .I0(ram16sdp_inst_132_dout[16]),
  .I1(ram16sdp_inst_140_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2041 (
  .O(mux_o_2041),
  .I0(ram16sdp_inst_148_dout[16]),
  .I1(ram16sdp_inst_156_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2042 (
  .O(mux_o_2042),
  .I0(ram16sdp_inst_164_dout[16]),
  .I1(ram16sdp_inst_172_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2043 (
  .O(mux_o_2043),
  .I0(ram16sdp_inst_180_dout[16]),
  .I1(ram16sdp_inst_188_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2044 (
  .O(mux_o_2044),
  .I0(ram16sdp_inst_196_dout[16]),
  .I1(ram16sdp_inst_204_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2045 (
  .O(mux_o_2045),
  .I0(ram16sdp_inst_212_dout[16]),
  .I1(ram16sdp_inst_220_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2046 (
  .O(mux_o_2046),
  .I0(ram16sdp_inst_228_dout[16]),
  .I1(ram16sdp_inst_236_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2047 (
  .O(mux_o_2047),
  .I0(ram16sdp_inst_244_dout[16]),
  .I1(ram16sdp_inst_252_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2048 (
  .O(mux_o_2048),
  .I0(ram16sdp_inst_260_dout[16]),
  .I1(ram16sdp_inst_268_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2049 (
  .O(mux_o_2049),
  .I0(ram16sdp_inst_276_dout[16]),
  .I1(ram16sdp_inst_284_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2050 (
  .O(mux_o_2050),
  .I0(ram16sdp_inst_292_dout[16]),
  .I1(ram16sdp_inst_300_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2051 (
  .O(mux_o_2051),
  .I0(ram16sdp_inst_308_dout[16]),
  .I1(ram16sdp_inst_316_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2052 (
  .O(mux_o_2052),
  .I0(ram16sdp_inst_324_dout[16]),
  .I1(ram16sdp_inst_332_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2053 (
  .O(mux_o_2053),
  .I0(ram16sdp_inst_340_dout[16]),
  .I1(ram16sdp_inst_348_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2054 (
  .O(mux_o_2054),
  .I0(ram16sdp_inst_356_dout[16]),
  .I1(ram16sdp_inst_364_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2055 (
  .O(mux_o_2055),
  .I0(ram16sdp_inst_372_dout[16]),
  .I1(ram16sdp_inst_380_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2056 (
  .O(mux_o_2056),
  .I0(ram16sdp_inst_388_dout[16]),
  .I1(ram16sdp_inst_396_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2057 (
  .O(mux_o_2057),
  .I0(ram16sdp_inst_404_dout[16]),
  .I1(ram16sdp_inst_412_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2058 (
  .O(mux_o_2058),
  .I0(ram16sdp_inst_420_dout[16]),
  .I1(ram16sdp_inst_428_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2059 (
  .O(mux_o_2059),
  .I0(ram16sdp_inst_436_dout[16]),
  .I1(ram16sdp_inst_444_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2060 (
  .O(mux_o_2060),
  .I0(ram16sdp_inst_452_dout[16]),
  .I1(ram16sdp_inst_460_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2061 (
  .O(mux_o_2061),
  .I0(ram16sdp_inst_468_dout[16]),
  .I1(ram16sdp_inst_476_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2062 (
  .O(mux_o_2062),
  .I0(ram16sdp_inst_484_dout[16]),
  .I1(ram16sdp_inst_492_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2063 (
  .O(mux_o_2063),
  .I0(ram16sdp_inst_500_dout[16]),
  .I1(ram16sdp_inst_508_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2064 (
  .O(mux_o_2064),
  .I0(ram16sdp_inst_516_dout[16]),
  .I1(ram16sdp_inst_524_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2065 (
  .O(mux_o_2065),
  .I0(ram16sdp_inst_532_dout[16]),
  .I1(ram16sdp_inst_540_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2066 (
  .O(mux_o_2066),
  .I0(ram16sdp_inst_548_dout[16]),
  .I1(ram16sdp_inst_556_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2067 (
  .O(mux_o_2067),
  .I0(ram16sdp_inst_564_dout[16]),
  .I1(ram16sdp_inst_572_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2068 (
  .O(mux_o_2068),
  .I0(ram16sdp_inst_580_dout[16]),
  .I1(ram16sdp_inst_588_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2069 (
  .O(mux_o_2069),
  .I0(ram16sdp_inst_596_dout[16]),
  .I1(ram16sdp_inst_604_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2070 (
  .O(mux_o_2070),
  .I0(ram16sdp_inst_612_dout[16]),
  .I1(ram16sdp_inst_620_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2071 (
  .O(mux_o_2071),
  .I0(ram16sdp_inst_628_dout[16]),
  .I1(ram16sdp_inst_636_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2072 (
  .O(mux_o_2072),
  .I0(ram16sdp_inst_644_dout[16]),
  .I1(ram16sdp_inst_652_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2073 (
  .O(mux_o_2073),
  .I0(ram16sdp_inst_660_dout[16]),
  .I1(ram16sdp_inst_668_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2074 (
  .O(mux_o_2074),
  .I0(ram16sdp_inst_676_dout[16]),
  .I1(ram16sdp_inst_684_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2075 (
  .O(mux_o_2075),
  .I0(ram16sdp_inst_692_dout[16]),
  .I1(ram16sdp_inst_700_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2076 (
  .O(mux_o_2076),
  .I0(ram16sdp_inst_708_dout[16]),
  .I1(ram16sdp_inst_716_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2077 (
  .O(mux_o_2077),
  .I0(ram16sdp_inst_724_dout[16]),
  .I1(ram16sdp_inst_732_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2078 (
  .O(mux_o_2078),
  .I0(ram16sdp_inst_740_dout[16]),
  .I1(ram16sdp_inst_748_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2079 (
  .O(mux_o_2079),
  .I0(ram16sdp_inst_756_dout[16]),
  .I1(ram16sdp_inst_764_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2080 (
  .O(mux_o_2080),
  .I0(ram16sdp_inst_772_dout[16]),
  .I1(ram16sdp_inst_780_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2081 (
  .O(mux_o_2081),
  .I0(ram16sdp_inst_788_dout[16]),
  .I1(ram16sdp_inst_796_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2082 (
  .O(mux_o_2082),
  .I0(ram16sdp_inst_804_dout[16]),
  .I1(ram16sdp_inst_812_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2083 (
  .O(mux_o_2083),
  .I0(ram16sdp_inst_820_dout[16]),
  .I1(ram16sdp_inst_828_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2084 (
  .O(mux_o_2084),
  .I0(ram16sdp_inst_836_dout[16]),
  .I1(ram16sdp_inst_844_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2085 (
  .O(mux_o_2085),
  .I0(ram16sdp_inst_852_dout[16]),
  .I1(ram16sdp_inst_860_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2086 (
  .O(mux_o_2086),
  .I0(ram16sdp_inst_868_dout[16]),
  .I1(ram16sdp_inst_876_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2087 (
  .O(mux_o_2087),
  .I0(ram16sdp_inst_884_dout[16]),
  .I1(ram16sdp_inst_892_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2088 (
  .O(mux_o_2088),
  .I0(ram16sdp_inst_900_dout[16]),
  .I1(ram16sdp_inst_908_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2089 (
  .O(mux_o_2089),
  .I0(ram16sdp_inst_916_dout[16]),
  .I1(ram16sdp_inst_924_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2090 (
  .O(mux_o_2090),
  .I0(ram16sdp_inst_932_dout[16]),
  .I1(ram16sdp_inst_940_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2091 (
  .O(mux_o_2091),
  .I0(ram16sdp_inst_948_dout[16]),
  .I1(ram16sdp_inst_956_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2092 (
  .O(mux_o_2092),
  .I0(ram16sdp_inst_964_dout[16]),
  .I1(ram16sdp_inst_972_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2093 (
  .O(mux_o_2093),
  .I0(ram16sdp_inst_980_dout[16]),
  .I1(ram16sdp_inst_988_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2094 (
  .O(mux_o_2094),
  .I0(ram16sdp_inst_996_dout[16]),
  .I1(ram16sdp_inst_1004_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2095 (
  .O(mux_o_2095),
  .I0(ram16sdp_inst_1012_dout[16]),
  .I1(ram16sdp_inst_1020_dout[16]),
  .S0(rad[4])
);
MUX2 mux_inst_2096 (
  .O(mux_o_2096),
  .I0(mux_o_2032),
  .I1(mux_o_2033),
  .S0(rad[5])
);
MUX2 mux_inst_2097 (
  .O(mux_o_2097),
  .I0(mux_o_2034),
  .I1(mux_o_2035),
  .S0(rad[5])
);
MUX2 mux_inst_2098 (
  .O(mux_o_2098),
  .I0(mux_o_2036),
  .I1(mux_o_2037),
  .S0(rad[5])
);
MUX2 mux_inst_2099 (
  .O(mux_o_2099),
  .I0(mux_o_2038),
  .I1(mux_o_2039),
  .S0(rad[5])
);
MUX2 mux_inst_2100 (
  .O(mux_o_2100),
  .I0(mux_o_2040),
  .I1(mux_o_2041),
  .S0(rad[5])
);
MUX2 mux_inst_2101 (
  .O(mux_o_2101),
  .I0(mux_o_2042),
  .I1(mux_o_2043),
  .S0(rad[5])
);
MUX2 mux_inst_2102 (
  .O(mux_o_2102),
  .I0(mux_o_2044),
  .I1(mux_o_2045),
  .S0(rad[5])
);
MUX2 mux_inst_2103 (
  .O(mux_o_2103),
  .I0(mux_o_2046),
  .I1(mux_o_2047),
  .S0(rad[5])
);
MUX2 mux_inst_2104 (
  .O(mux_o_2104),
  .I0(mux_o_2048),
  .I1(mux_o_2049),
  .S0(rad[5])
);
MUX2 mux_inst_2105 (
  .O(mux_o_2105),
  .I0(mux_o_2050),
  .I1(mux_o_2051),
  .S0(rad[5])
);
MUX2 mux_inst_2106 (
  .O(mux_o_2106),
  .I0(mux_o_2052),
  .I1(mux_o_2053),
  .S0(rad[5])
);
MUX2 mux_inst_2107 (
  .O(mux_o_2107),
  .I0(mux_o_2054),
  .I1(mux_o_2055),
  .S0(rad[5])
);
MUX2 mux_inst_2108 (
  .O(mux_o_2108),
  .I0(mux_o_2056),
  .I1(mux_o_2057),
  .S0(rad[5])
);
MUX2 mux_inst_2109 (
  .O(mux_o_2109),
  .I0(mux_o_2058),
  .I1(mux_o_2059),
  .S0(rad[5])
);
MUX2 mux_inst_2110 (
  .O(mux_o_2110),
  .I0(mux_o_2060),
  .I1(mux_o_2061),
  .S0(rad[5])
);
MUX2 mux_inst_2111 (
  .O(mux_o_2111),
  .I0(mux_o_2062),
  .I1(mux_o_2063),
  .S0(rad[5])
);
MUX2 mux_inst_2112 (
  .O(mux_o_2112),
  .I0(mux_o_2064),
  .I1(mux_o_2065),
  .S0(rad[5])
);
MUX2 mux_inst_2113 (
  .O(mux_o_2113),
  .I0(mux_o_2066),
  .I1(mux_o_2067),
  .S0(rad[5])
);
MUX2 mux_inst_2114 (
  .O(mux_o_2114),
  .I0(mux_o_2068),
  .I1(mux_o_2069),
  .S0(rad[5])
);
MUX2 mux_inst_2115 (
  .O(mux_o_2115),
  .I0(mux_o_2070),
  .I1(mux_o_2071),
  .S0(rad[5])
);
MUX2 mux_inst_2116 (
  .O(mux_o_2116),
  .I0(mux_o_2072),
  .I1(mux_o_2073),
  .S0(rad[5])
);
MUX2 mux_inst_2117 (
  .O(mux_o_2117),
  .I0(mux_o_2074),
  .I1(mux_o_2075),
  .S0(rad[5])
);
MUX2 mux_inst_2118 (
  .O(mux_o_2118),
  .I0(mux_o_2076),
  .I1(mux_o_2077),
  .S0(rad[5])
);
MUX2 mux_inst_2119 (
  .O(mux_o_2119),
  .I0(mux_o_2078),
  .I1(mux_o_2079),
  .S0(rad[5])
);
MUX2 mux_inst_2120 (
  .O(mux_o_2120),
  .I0(mux_o_2080),
  .I1(mux_o_2081),
  .S0(rad[5])
);
MUX2 mux_inst_2121 (
  .O(mux_o_2121),
  .I0(mux_o_2082),
  .I1(mux_o_2083),
  .S0(rad[5])
);
MUX2 mux_inst_2122 (
  .O(mux_o_2122),
  .I0(mux_o_2084),
  .I1(mux_o_2085),
  .S0(rad[5])
);
MUX2 mux_inst_2123 (
  .O(mux_o_2123),
  .I0(mux_o_2086),
  .I1(mux_o_2087),
  .S0(rad[5])
);
MUX2 mux_inst_2124 (
  .O(mux_o_2124),
  .I0(mux_o_2088),
  .I1(mux_o_2089),
  .S0(rad[5])
);
MUX2 mux_inst_2125 (
  .O(mux_o_2125),
  .I0(mux_o_2090),
  .I1(mux_o_2091),
  .S0(rad[5])
);
MUX2 mux_inst_2126 (
  .O(mux_o_2126),
  .I0(mux_o_2092),
  .I1(mux_o_2093),
  .S0(rad[5])
);
MUX2 mux_inst_2127 (
  .O(mux_o_2127),
  .I0(mux_o_2094),
  .I1(mux_o_2095),
  .S0(rad[5])
);
MUX2 mux_inst_2128 (
  .O(mux_o_2128),
  .I0(mux_o_2096),
  .I1(mux_o_2097),
  .S0(rad[6])
);
MUX2 mux_inst_2129 (
  .O(mux_o_2129),
  .I0(mux_o_2098),
  .I1(mux_o_2099),
  .S0(rad[6])
);
MUX2 mux_inst_2130 (
  .O(mux_o_2130),
  .I0(mux_o_2100),
  .I1(mux_o_2101),
  .S0(rad[6])
);
MUX2 mux_inst_2131 (
  .O(mux_o_2131),
  .I0(mux_o_2102),
  .I1(mux_o_2103),
  .S0(rad[6])
);
MUX2 mux_inst_2132 (
  .O(mux_o_2132),
  .I0(mux_o_2104),
  .I1(mux_o_2105),
  .S0(rad[6])
);
MUX2 mux_inst_2133 (
  .O(mux_o_2133),
  .I0(mux_o_2106),
  .I1(mux_o_2107),
  .S0(rad[6])
);
MUX2 mux_inst_2134 (
  .O(mux_o_2134),
  .I0(mux_o_2108),
  .I1(mux_o_2109),
  .S0(rad[6])
);
MUX2 mux_inst_2135 (
  .O(mux_o_2135),
  .I0(mux_o_2110),
  .I1(mux_o_2111),
  .S0(rad[6])
);
MUX2 mux_inst_2136 (
  .O(mux_o_2136),
  .I0(mux_o_2112),
  .I1(mux_o_2113),
  .S0(rad[6])
);
MUX2 mux_inst_2137 (
  .O(mux_o_2137),
  .I0(mux_o_2114),
  .I1(mux_o_2115),
  .S0(rad[6])
);
MUX2 mux_inst_2138 (
  .O(mux_o_2138),
  .I0(mux_o_2116),
  .I1(mux_o_2117),
  .S0(rad[6])
);
MUX2 mux_inst_2139 (
  .O(mux_o_2139),
  .I0(mux_o_2118),
  .I1(mux_o_2119),
  .S0(rad[6])
);
MUX2 mux_inst_2140 (
  .O(mux_o_2140),
  .I0(mux_o_2120),
  .I1(mux_o_2121),
  .S0(rad[6])
);
MUX2 mux_inst_2141 (
  .O(mux_o_2141),
  .I0(mux_o_2122),
  .I1(mux_o_2123),
  .S0(rad[6])
);
MUX2 mux_inst_2142 (
  .O(mux_o_2142),
  .I0(mux_o_2124),
  .I1(mux_o_2125),
  .S0(rad[6])
);
MUX2 mux_inst_2143 (
  .O(mux_o_2143),
  .I0(mux_o_2126),
  .I1(mux_o_2127),
  .S0(rad[6])
);
MUX2 mux_inst_2144 (
  .O(mux_o_2144),
  .I0(mux_o_2128),
  .I1(mux_o_2129),
  .S0(rad[7])
);
MUX2 mux_inst_2145 (
  .O(mux_o_2145),
  .I0(mux_o_2130),
  .I1(mux_o_2131),
  .S0(rad[7])
);
MUX2 mux_inst_2146 (
  .O(mux_o_2146),
  .I0(mux_o_2132),
  .I1(mux_o_2133),
  .S0(rad[7])
);
MUX2 mux_inst_2147 (
  .O(mux_o_2147),
  .I0(mux_o_2134),
  .I1(mux_o_2135),
  .S0(rad[7])
);
MUX2 mux_inst_2148 (
  .O(mux_o_2148),
  .I0(mux_o_2136),
  .I1(mux_o_2137),
  .S0(rad[7])
);
MUX2 mux_inst_2149 (
  .O(mux_o_2149),
  .I0(mux_o_2138),
  .I1(mux_o_2139),
  .S0(rad[7])
);
MUX2 mux_inst_2150 (
  .O(mux_o_2150),
  .I0(mux_o_2140),
  .I1(mux_o_2141),
  .S0(rad[7])
);
MUX2 mux_inst_2151 (
  .O(mux_o_2151),
  .I0(mux_o_2142),
  .I1(mux_o_2143),
  .S0(rad[7])
);
MUX2 mux_inst_2152 (
  .O(mux_o_2152),
  .I0(mux_o_2144),
  .I1(mux_o_2145),
  .S0(rad[8])
);
MUX2 mux_inst_2153 (
  .O(mux_o_2153),
  .I0(mux_o_2146),
  .I1(mux_o_2147),
  .S0(rad[8])
);
MUX2 mux_inst_2154 (
  .O(mux_o_2154),
  .I0(mux_o_2148),
  .I1(mux_o_2149),
  .S0(rad[8])
);
MUX2 mux_inst_2155 (
  .O(mux_o_2155),
  .I0(mux_o_2150),
  .I1(mux_o_2151),
  .S0(rad[8])
);
MUX2 mux_inst_2156 (
  .O(mux_o_2156),
  .I0(mux_o_2152),
  .I1(mux_o_2153),
  .S0(rad[9])
);
MUX2 mux_inst_2157 (
  .O(mux_o_2157),
  .I0(mux_o_2154),
  .I1(mux_o_2155),
  .S0(rad[9])
);
MUX2 mux_inst_2158 (
  .O(dout[16]),
  .I0(mux_o_2156),
  .I1(mux_o_2157),
  .S0(rad[10])
);
MUX2 mux_inst_2159 (
  .O(mux_o_2159),
  .I0(ram16sdp_inst_4_dout[17]),
  .I1(ram16sdp_inst_12_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2160 (
  .O(mux_o_2160),
  .I0(ram16sdp_inst_20_dout[17]),
  .I1(ram16sdp_inst_28_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2161 (
  .O(mux_o_2161),
  .I0(ram16sdp_inst_36_dout[17]),
  .I1(ram16sdp_inst_44_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2162 (
  .O(mux_o_2162),
  .I0(ram16sdp_inst_52_dout[17]),
  .I1(ram16sdp_inst_60_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2163 (
  .O(mux_o_2163),
  .I0(ram16sdp_inst_68_dout[17]),
  .I1(ram16sdp_inst_76_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2164 (
  .O(mux_o_2164),
  .I0(ram16sdp_inst_84_dout[17]),
  .I1(ram16sdp_inst_92_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2165 (
  .O(mux_o_2165),
  .I0(ram16sdp_inst_100_dout[17]),
  .I1(ram16sdp_inst_108_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2166 (
  .O(mux_o_2166),
  .I0(ram16sdp_inst_116_dout[17]),
  .I1(ram16sdp_inst_124_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2167 (
  .O(mux_o_2167),
  .I0(ram16sdp_inst_132_dout[17]),
  .I1(ram16sdp_inst_140_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2168 (
  .O(mux_o_2168),
  .I0(ram16sdp_inst_148_dout[17]),
  .I1(ram16sdp_inst_156_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2169 (
  .O(mux_o_2169),
  .I0(ram16sdp_inst_164_dout[17]),
  .I1(ram16sdp_inst_172_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2170 (
  .O(mux_o_2170),
  .I0(ram16sdp_inst_180_dout[17]),
  .I1(ram16sdp_inst_188_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2171 (
  .O(mux_o_2171),
  .I0(ram16sdp_inst_196_dout[17]),
  .I1(ram16sdp_inst_204_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2172 (
  .O(mux_o_2172),
  .I0(ram16sdp_inst_212_dout[17]),
  .I1(ram16sdp_inst_220_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2173 (
  .O(mux_o_2173),
  .I0(ram16sdp_inst_228_dout[17]),
  .I1(ram16sdp_inst_236_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2174 (
  .O(mux_o_2174),
  .I0(ram16sdp_inst_244_dout[17]),
  .I1(ram16sdp_inst_252_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2175 (
  .O(mux_o_2175),
  .I0(ram16sdp_inst_260_dout[17]),
  .I1(ram16sdp_inst_268_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2176 (
  .O(mux_o_2176),
  .I0(ram16sdp_inst_276_dout[17]),
  .I1(ram16sdp_inst_284_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2177 (
  .O(mux_o_2177),
  .I0(ram16sdp_inst_292_dout[17]),
  .I1(ram16sdp_inst_300_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2178 (
  .O(mux_o_2178),
  .I0(ram16sdp_inst_308_dout[17]),
  .I1(ram16sdp_inst_316_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2179 (
  .O(mux_o_2179),
  .I0(ram16sdp_inst_324_dout[17]),
  .I1(ram16sdp_inst_332_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2180 (
  .O(mux_o_2180),
  .I0(ram16sdp_inst_340_dout[17]),
  .I1(ram16sdp_inst_348_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2181 (
  .O(mux_o_2181),
  .I0(ram16sdp_inst_356_dout[17]),
  .I1(ram16sdp_inst_364_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2182 (
  .O(mux_o_2182),
  .I0(ram16sdp_inst_372_dout[17]),
  .I1(ram16sdp_inst_380_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2183 (
  .O(mux_o_2183),
  .I0(ram16sdp_inst_388_dout[17]),
  .I1(ram16sdp_inst_396_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2184 (
  .O(mux_o_2184),
  .I0(ram16sdp_inst_404_dout[17]),
  .I1(ram16sdp_inst_412_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2185 (
  .O(mux_o_2185),
  .I0(ram16sdp_inst_420_dout[17]),
  .I1(ram16sdp_inst_428_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2186 (
  .O(mux_o_2186),
  .I0(ram16sdp_inst_436_dout[17]),
  .I1(ram16sdp_inst_444_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2187 (
  .O(mux_o_2187),
  .I0(ram16sdp_inst_452_dout[17]),
  .I1(ram16sdp_inst_460_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2188 (
  .O(mux_o_2188),
  .I0(ram16sdp_inst_468_dout[17]),
  .I1(ram16sdp_inst_476_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2189 (
  .O(mux_o_2189),
  .I0(ram16sdp_inst_484_dout[17]),
  .I1(ram16sdp_inst_492_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2190 (
  .O(mux_o_2190),
  .I0(ram16sdp_inst_500_dout[17]),
  .I1(ram16sdp_inst_508_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2191 (
  .O(mux_o_2191),
  .I0(ram16sdp_inst_516_dout[17]),
  .I1(ram16sdp_inst_524_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2192 (
  .O(mux_o_2192),
  .I0(ram16sdp_inst_532_dout[17]),
  .I1(ram16sdp_inst_540_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2193 (
  .O(mux_o_2193),
  .I0(ram16sdp_inst_548_dout[17]),
  .I1(ram16sdp_inst_556_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2194 (
  .O(mux_o_2194),
  .I0(ram16sdp_inst_564_dout[17]),
  .I1(ram16sdp_inst_572_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2195 (
  .O(mux_o_2195),
  .I0(ram16sdp_inst_580_dout[17]),
  .I1(ram16sdp_inst_588_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2196 (
  .O(mux_o_2196),
  .I0(ram16sdp_inst_596_dout[17]),
  .I1(ram16sdp_inst_604_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2197 (
  .O(mux_o_2197),
  .I0(ram16sdp_inst_612_dout[17]),
  .I1(ram16sdp_inst_620_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2198 (
  .O(mux_o_2198),
  .I0(ram16sdp_inst_628_dout[17]),
  .I1(ram16sdp_inst_636_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2199 (
  .O(mux_o_2199),
  .I0(ram16sdp_inst_644_dout[17]),
  .I1(ram16sdp_inst_652_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2200 (
  .O(mux_o_2200),
  .I0(ram16sdp_inst_660_dout[17]),
  .I1(ram16sdp_inst_668_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2201 (
  .O(mux_o_2201),
  .I0(ram16sdp_inst_676_dout[17]),
  .I1(ram16sdp_inst_684_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2202 (
  .O(mux_o_2202),
  .I0(ram16sdp_inst_692_dout[17]),
  .I1(ram16sdp_inst_700_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2203 (
  .O(mux_o_2203),
  .I0(ram16sdp_inst_708_dout[17]),
  .I1(ram16sdp_inst_716_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2204 (
  .O(mux_o_2204),
  .I0(ram16sdp_inst_724_dout[17]),
  .I1(ram16sdp_inst_732_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2205 (
  .O(mux_o_2205),
  .I0(ram16sdp_inst_740_dout[17]),
  .I1(ram16sdp_inst_748_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2206 (
  .O(mux_o_2206),
  .I0(ram16sdp_inst_756_dout[17]),
  .I1(ram16sdp_inst_764_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2207 (
  .O(mux_o_2207),
  .I0(ram16sdp_inst_772_dout[17]),
  .I1(ram16sdp_inst_780_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2208 (
  .O(mux_o_2208),
  .I0(ram16sdp_inst_788_dout[17]),
  .I1(ram16sdp_inst_796_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2209 (
  .O(mux_o_2209),
  .I0(ram16sdp_inst_804_dout[17]),
  .I1(ram16sdp_inst_812_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2210 (
  .O(mux_o_2210),
  .I0(ram16sdp_inst_820_dout[17]),
  .I1(ram16sdp_inst_828_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2211 (
  .O(mux_o_2211),
  .I0(ram16sdp_inst_836_dout[17]),
  .I1(ram16sdp_inst_844_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2212 (
  .O(mux_o_2212),
  .I0(ram16sdp_inst_852_dout[17]),
  .I1(ram16sdp_inst_860_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2213 (
  .O(mux_o_2213),
  .I0(ram16sdp_inst_868_dout[17]),
  .I1(ram16sdp_inst_876_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2214 (
  .O(mux_o_2214),
  .I0(ram16sdp_inst_884_dout[17]),
  .I1(ram16sdp_inst_892_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2215 (
  .O(mux_o_2215),
  .I0(ram16sdp_inst_900_dout[17]),
  .I1(ram16sdp_inst_908_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2216 (
  .O(mux_o_2216),
  .I0(ram16sdp_inst_916_dout[17]),
  .I1(ram16sdp_inst_924_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2217 (
  .O(mux_o_2217),
  .I0(ram16sdp_inst_932_dout[17]),
  .I1(ram16sdp_inst_940_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2218 (
  .O(mux_o_2218),
  .I0(ram16sdp_inst_948_dout[17]),
  .I1(ram16sdp_inst_956_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2219 (
  .O(mux_o_2219),
  .I0(ram16sdp_inst_964_dout[17]),
  .I1(ram16sdp_inst_972_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2220 (
  .O(mux_o_2220),
  .I0(ram16sdp_inst_980_dout[17]),
  .I1(ram16sdp_inst_988_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2221 (
  .O(mux_o_2221),
  .I0(ram16sdp_inst_996_dout[17]),
  .I1(ram16sdp_inst_1004_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2222 (
  .O(mux_o_2222),
  .I0(ram16sdp_inst_1012_dout[17]),
  .I1(ram16sdp_inst_1020_dout[17]),
  .S0(rad[4])
);
MUX2 mux_inst_2223 (
  .O(mux_o_2223),
  .I0(mux_o_2159),
  .I1(mux_o_2160),
  .S0(rad[5])
);
MUX2 mux_inst_2224 (
  .O(mux_o_2224),
  .I0(mux_o_2161),
  .I1(mux_o_2162),
  .S0(rad[5])
);
MUX2 mux_inst_2225 (
  .O(mux_o_2225),
  .I0(mux_o_2163),
  .I1(mux_o_2164),
  .S0(rad[5])
);
MUX2 mux_inst_2226 (
  .O(mux_o_2226),
  .I0(mux_o_2165),
  .I1(mux_o_2166),
  .S0(rad[5])
);
MUX2 mux_inst_2227 (
  .O(mux_o_2227),
  .I0(mux_o_2167),
  .I1(mux_o_2168),
  .S0(rad[5])
);
MUX2 mux_inst_2228 (
  .O(mux_o_2228),
  .I0(mux_o_2169),
  .I1(mux_o_2170),
  .S0(rad[5])
);
MUX2 mux_inst_2229 (
  .O(mux_o_2229),
  .I0(mux_o_2171),
  .I1(mux_o_2172),
  .S0(rad[5])
);
MUX2 mux_inst_2230 (
  .O(mux_o_2230),
  .I0(mux_o_2173),
  .I1(mux_o_2174),
  .S0(rad[5])
);
MUX2 mux_inst_2231 (
  .O(mux_o_2231),
  .I0(mux_o_2175),
  .I1(mux_o_2176),
  .S0(rad[5])
);
MUX2 mux_inst_2232 (
  .O(mux_o_2232),
  .I0(mux_o_2177),
  .I1(mux_o_2178),
  .S0(rad[5])
);
MUX2 mux_inst_2233 (
  .O(mux_o_2233),
  .I0(mux_o_2179),
  .I1(mux_o_2180),
  .S0(rad[5])
);
MUX2 mux_inst_2234 (
  .O(mux_o_2234),
  .I0(mux_o_2181),
  .I1(mux_o_2182),
  .S0(rad[5])
);
MUX2 mux_inst_2235 (
  .O(mux_o_2235),
  .I0(mux_o_2183),
  .I1(mux_o_2184),
  .S0(rad[5])
);
MUX2 mux_inst_2236 (
  .O(mux_o_2236),
  .I0(mux_o_2185),
  .I1(mux_o_2186),
  .S0(rad[5])
);
MUX2 mux_inst_2237 (
  .O(mux_o_2237),
  .I0(mux_o_2187),
  .I1(mux_o_2188),
  .S0(rad[5])
);
MUX2 mux_inst_2238 (
  .O(mux_o_2238),
  .I0(mux_o_2189),
  .I1(mux_o_2190),
  .S0(rad[5])
);
MUX2 mux_inst_2239 (
  .O(mux_o_2239),
  .I0(mux_o_2191),
  .I1(mux_o_2192),
  .S0(rad[5])
);
MUX2 mux_inst_2240 (
  .O(mux_o_2240),
  .I0(mux_o_2193),
  .I1(mux_o_2194),
  .S0(rad[5])
);
MUX2 mux_inst_2241 (
  .O(mux_o_2241),
  .I0(mux_o_2195),
  .I1(mux_o_2196),
  .S0(rad[5])
);
MUX2 mux_inst_2242 (
  .O(mux_o_2242),
  .I0(mux_o_2197),
  .I1(mux_o_2198),
  .S0(rad[5])
);
MUX2 mux_inst_2243 (
  .O(mux_o_2243),
  .I0(mux_o_2199),
  .I1(mux_o_2200),
  .S0(rad[5])
);
MUX2 mux_inst_2244 (
  .O(mux_o_2244),
  .I0(mux_o_2201),
  .I1(mux_o_2202),
  .S0(rad[5])
);
MUX2 mux_inst_2245 (
  .O(mux_o_2245),
  .I0(mux_o_2203),
  .I1(mux_o_2204),
  .S0(rad[5])
);
MUX2 mux_inst_2246 (
  .O(mux_o_2246),
  .I0(mux_o_2205),
  .I1(mux_o_2206),
  .S0(rad[5])
);
MUX2 mux_inst_2247 (
  .O(mux_o_2247),
  .I0(mux_o_2207),
  .I1(mux_o_2208),
  .S0(rad[5])
);
MUX2 mux_inst_2248 (
  .O(mux_o_2248),
  .I0(mux_o_2209),
  .I1(mux_o_2210),
  .S0(rad[5])
);
MUX2 mux_inst_2249 (
  .O(mux_o_2249),
  .I0(mux_o_2211),
  .I1(mux_o_2212),
  .S0(rad[5])
);
MUX2 mux_inst_2250 (
  .O(mux_o_2250),
  .I0(mux_o_2213),
  .I1(mux_o_2214),
  .S0(rad[5])
);
MUX2 mux_inst_2251 (
  .O(mux_o_2251),
  .I0(mux_o_2215),
  .I1(mux_o_2216),
  .S0(rad[5])
);
MUX2 mux_inst_2252 (
  .O(mux_o_2252),
  .I0(mux_o_2217),
  .I1(mux_o_2218),
  .S0(rad[5])
);
MUX2 mux_inst_2253 (
  .O(mux_o_2253),
  .I0(mux_o_2219),
  .I1(mux_o_2220),
  .S0(rad[5])
);
MUX2 mux_inst_2254 (
  .O(mux_o_2254),
  .I0(mux_o_2221),
  .I1(mux_o_2222),
  .S0(rad[5])
);
MUX2 mux_inst_2255 (
  .O(mux_o_2255),
  .I0(mux_o_2223),
  .I1(mux_o_2224),
  .S0(rad[6])
);
MUX2 mux_inst_2256 (
  .O(mux_o_2256),
  .I0(mux_o_2225),
  .I1(mux_o_2226),
  .S0(rad[6])
);
MUX2 mux_inst_2257 (
  .O(mux_o_2257),
  .I0(mux_o_2227),
  .I1(mux_o_2228),
  .S0(rad[6])
);
MUX2 mux_inst_2258 (
  .O(mux_o_2258),
  .I0(mux_o_2229),
  .I1(mux_o_2230),
  .S0(rad[6])
);
MUX2 mux_inst_2259 (
  .O(mux_o_2259),
  .I0(mux_o_2231),
  .I1(mux_o_2232),
  .S0(rad[6])
);
MUX2 mux_inst_2260 (
  .O(mux_o_2260),
  .I0(mux_o_2233),
  .I1(mux_o_2234),
  .S0(rad[6])
);
MUX2 mux_inst_2261 (
  .O(mux_o_2261),
  .I0(mux_o_2235),
  .I1(mux_o_2236),
  .S0(rad[6])
);
MUX2 mux_inst_2262 (
  .O(mux_o_2262),
  .I0(mux_o_2237),
  .I1(mux_o_2238),
  .S0(rad[6])
);
MUX2 mux_inst_2263 (
  .O(mux_o_2263),
  .I0(mux_o_2239),
  .I1(mux_o_2240),
  .S0(rad[6])
);
MUX2 mux_inst_2264 (
  .O(mux_o_2264),
  .I0(mux_o_2241),
  .I1(mux_o_2242),
  .S0(rad[6])
);
MUX2 mux_inst_2265 (
  .O(mux_o_2265),
  .I0(mux_o_2243),
  .I1(mux_o_2244),
  .S0(rad[6])
);
MUX2 mux_inst_2266 (
  .O(mux_o_2266),
  .I0(mux_o_2245),
  .I1(mux_o_2246),
  .S0(rad[6])
);
MUX2 mux_inst_2267 (
  .O(mux_o_2267),
  .I0(mux_o_2247),
  .I1(mux_o_2248),
  .S0(rad[6])
);
MUX2 mux_inst_2268 (
  .O(mux_o_2268),
  .I0(mux_o_2249),
  .I1(mux_o_2250),
  .S0(rad[6])
);
MUX2 mux_inst_2269 (
  .O(mux_o_2269),
  .I0(mux_o_2251),
  .I1(mux_o_2252),
  .S0(rad[6])
);
MUX2 mux_inst_2270 (
  .O(mux_o_2270),
  .I0(mux_o_2253),
  .I1(mux_o_2254),
  .S0(rad[6])
);
MUX2 mux_inst_2271 (
  .O(mux_o_2271),
  .I0(mux_o_2255),
  .I1(mux_o_2256),
  .S0(rad[7])
);
MUX2 mux_inst_2272 (
  .O(mux_o_2272),
  .I0(mux_o_2257),
  .I1(mux_o_2258),
  .S0(rad[7])
);
MUX2 mux_inst_2273 (
  .O(mux_o_2273),
  .I0(mux_o_2259),
  .I1(mux_o_2260),
  .S0(rad[7])
);
MUX2 mux_inst_2274 (
  .O(mux_o_2274),
  .I0(mux_o_2261),
  .I1(mux_o_2262),
  .S0(rad[7])
);
MUX2 mux_inst_2275 (
  .O(mux_o_2275),
  .I0(mux_o_2263),
  .I1(mux_o_2264),
  .S0(rad[7])
);
MUX2 mux_inst_2276 (
  .O(mux_o_2276),
  .I0(mux_o_2265),
  .I1(mux_o_2266),
  .S0(rad[7])
);
MUX2 mux_inst_2277 (
  .O(mux_o_2277),
  .I0(mux_o_2267),
  .I1(mux_o_2268),
  .S0(rad[7])
);
MUX2 mux_inst_2278 (
  .O(mux_o_2278),
  .I0(mux_o_2269),
  .I1(mux_o_2270),
  .S0(rad[7])
);
MUX2 mux_inst_2279 (
  .O(mux_o_2279),
  .I0(mux_o_2271),
  .I1(mux_o_2272),
  .S0(rad[8])
);
MUX2 mux_inst_2280 (
  .O(mux_o_2280),
  .I0(mux_o_2273),
  .I1(mux_o_2274),
  .S0(rad[8])
);
MUX2 mux_inst_2281 (
  .O(mux_o_2281),
  .I0(mux_o_2275),
  .I1(mux_o_2276),
  .S0(rad[8])
);
MUX2 mux_inst_2282 (
  .O(mux_o_2282),
  .I0(mux_o_2277),
  .I1(mux_o_2278),
  .S0(rad[8])
);
MUX2 mux_inst_2283 (
  .O(mux_o_2283),
  .I0(mux_o_2279),
  .I1(mux_o_2280),
  .S0(rad[9])
);
MUX2 mux_inst_2284 (
  .O(mux_o_2284),
  .I0(mux_o_2281),
  .I1(mux_o_2282),
  .S0(rad[9])
);
MUX2 mux_inst_2285 (
  .O(dout[17]),
  .I0(mux_o_2283),
  .I1(mux_o_2284),
  .S0(rad[10])
);
MUX2 mux_inst_2286 (
  .O(mux_o_2286),
  .I0(ram16sdp_inst_4_dout[18]),
  .I1(ram16sdp_inst_12_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2287 (
  .O(mux_o_2287),
  .I0(ram16sdp_inst_20_dout[18]),
  .I1(ram16sdp_inst_28_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2288 (
  .O(mux_o_2288),
  .I0(ram16sdp_inst_36_dout[18]),
  .I1(ram16sdp_inst_44_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2289 (
  .O(mux_o_2289),
  .I0(ram16sdp_inst_52_dout[18]),
  .I1(ram16sdp_inst_60_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2290 (
  .O(mux_o_2290),
  .I0(ram16sdp_inst_68_dout[18]),
  .I1(ram16sdp_inst_76_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2291 (
  .O(mux_o_2291),
  .I0(ram16sdp_inst_84_dout[18]),
  .I1(ram16sdp_inst_92_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2292 (
  .O(mux_o_2292),
  .I0(ram16sdp_inst_100_dout[18]),
  .I1(ram16sdp_inst_108_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2293 (
  .O(mux_o_2293),
  .I0(ram16sdp_inst_116_dout[18]),
  .I1(ram16sdp_inst_124_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2294 (
  .O(mux_o_2294),
  .I0(ram16sdp_inst_132_dout[18]),
  .I1(ram16sdp_inst_140_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2295 (
  .O(mux_o_2295),
  .I0(ram16sdp_inst_148_dout[18]),
  .I1(ram16sdp_inst_156_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2296 (
  .O(mux_o_2296),
  .I0(ram16sdp_inst_164_dout[18]),
  .I1(ram16sdp_inst_172_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2297 (
  .O(mux_o_2297),
  .I0(ram16sdp_inst_180_dout[18]),
  .I1(ram16sdp_inst_188_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2298 (
  .O(mux_o_2298),
  .I0(ram16sdp_inst_196_dout[18]),
  .I1(ram16sdp_inst_204_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2299 (
  .O(mux_o_2299),
  .I0(ram16sdp_inst_212_dout[18]),
  .I1(ram16sdp_inst_220_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2300 (
  .O(mux_o_2300),
  .I0(ram16sdp_inst_228_dout[18]),
  .I1(ram16sdp_inst_236_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2301 (
  .O(mux_o_2301),
  .I0(ram16sdp_inst_244_dout[18]),
  .I1(ram16sdp_inst_252_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2302 (
  .O(mux_o_2302),
  .I0(ram16sdp_inst_260_dout[18]),
  .I1(ram16sdp_inst_268_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2303 (
  .O(mux_o_2303),
  .I0(ram16sdp_inst_276_dout[18]),
  .I1(ram16sdp_inst_284_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2304 (
  .O(mux_o_2304),
  .I0(ram16sdp_inst_292_dout[18]),
  .I1(ram16sdp_inst_300_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2305 (
  .O(mux_o_2305),
  .I0(ram16sdp_inst_308_dout[18]),
  .I1(ram16sdp_inst_316_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2306 (
  .O(mux_o_2306),
  .I0(ram16sdp_inst_324_dout[18]),
  .I1(ram16sdp_inst_332_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2307 (
  .O(mux_o_2307),
  .I0(ram16sdp_inst_340_dout[18]),
  .I1(ram16sdp_inst_348_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2308 (
  .O(mux_o_2308),
  .I0(ram16sdp_inst_356_dout[18]),
  .I1(ram16sdp_inst_364_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2309 (
  .O(mux_o_2309),
  .I0(ram16sdp_inst_372_dout[18]),
  .I1(ram16sdp_inst_380_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2310 (
  .O(mux_o_2310),
  .I0(ram16sdp_inst_388_dout[18]),
  .I1(ram16sdp_inst_396_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2311 (
  .O(mux_o_2311),
  .I0(ram16sdp_inst_404_dout[18]),
  .I1(ram16sdp_inst_412_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2312 (
  .O(mux_o_2312),
  .I0(ram16sdp_inst_420_dout[18]),
  .I1(ram16sdp_inst_428_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2313 (
  .O(mux_o_2313),
  .I0(ram16sdp_inst_436_dout[18]),
  .I1(ram16sdp_inst_444_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2314 (
  .O(mux_o_2314),
  .I0(ram16sdp_inst_452_dout[18]),
  .I1(ram16sdp_inst_460_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2315 (
  .O(mux_o_2315),
  .I0(ram16sdp_inst_468_dout[18]),
  .I1(ram16sdp_inst_476_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2316 (
  .O(mux_o_2316),
  .I0(ram16sdp_inst_484_dout[18]),
  .I1(ram16sdp_inst_492_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2317 (
  .O(mux_o_2317),
  .I0(ram16sdp_inst_500_dout[18]),
  .I1(ram16sdp_inst_508_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2318 (
  .O(mux_o_2318),
  .I0(ram16sdp_inst_516_dout[18]),
  .I1(ram16sdp_inst_524_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2319 (
  .O(mux_o_2319),
  .I0(ram16sdp_inst_532_dout[18]),
  .I1(ram16sdp_inst_540_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2320 (
  .O(mux_o_2320),
  .I0(ram16sdp_inst_548_dout[18]),
  .I1(ram16sdp_inst_556_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2321 (
  .O(mux_o_2321),
  .I0(ram16sdp_inst_564_dout[18]),
  .I1(ram16sdp_inst_572_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2322 (
  .O(mux_o_2322),
  .I0(ram16sdp_inst_580_dout[18]),
  .I1(ram16sdp_inst_588_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2323 (
  .O(mux_o_2323),
  .I0(ram16sdp_inst_596_dout[18]),
  .I1(ram16sdp_inst_604_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2324 (
  .O(mux_o_2324),
  .I0(ram16sdp_inst_612_dout[18]),
  .I1(ram16sdp_inst_620_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2325 (
  .O(mux_o_2325),
  .I0(ram16sdp_inst_628_dout[18]),
  .I1(ram16sdp_inst_636_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2326 (
  .O(mux_o_2326),
  .I0(ram16sdp_inst_644_dout[18]),
  .I1(ram16sdp_inst_652_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2327 (
  .O(mux_o_2327),
  .I0(ram16sdp_inst_660_dout[18]),
  .I1(ram16sdp_inst_668_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2328 (
  .O(mux_o_2328),
  .I0(ram16sdp_inst_676_dout[18]),
  .I1(ram16sdp_inst_684_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2329 (
  .O(mux_o_2329),
  .I0(ram16sdp_inst_692_dout[18]),
  .I1(ram16sdp_inst_700_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2330 (
  .O(mux_o_2330),
  .I0(ram16sdp_inst_708_dout[18]),
  .I1(ram16sdp_inst_716_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2331 (
  .O(mux_o_2331),
  .I0(ram16sdp_inst_724_dout[18]),
  .I1(ram16sdp_inst_732_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2332 (
  .O(mux_o_2332),
  .I0(ram16sdp_inst_740_dout[18]),
  .I1(ram16sdp_inst_748_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2333 (
  .O(mux_o_2333),
  .I0(ram16sdp_inst_756_dout[18]),
  .I1(ram16sdp_inst_764_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2334 (
  .O(mux_o_2334),
  .I0(ram16sdp_inst_772_dout[18]),
  .I1(ram16sdp_inst_780_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2335 (
  .O(mux_o_2335),
  .I0(ram16sdp_inst_788_dout[18]),
  .I1(ram16sdp_inst_796_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2336 (
  .O(mux_o_2336),
  .I0(ram16sdp_inst_804_dout[18]),
  .I1(ram16sdp_inst_812_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2337 (
  .O(mux_o_2337),
  .I0(ram16sdp_inst_820_dout[18]),
  .I1(ram16sdp_inst_828_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2338 (
  .O(mux_o_2338),
  .I0(ram16sdp_inst_836_dout[18]),
  .I1(ram16sdp_inst_844_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2339 (
  .O(mux_o_2339),
  .I0(ram16sdp_inst_852_dout[18]),
  .I1(ram16sdp_inst_860_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2340 (
  .O(mux_o_2340),
  .I0(ram16sdp_inst_868_dout[18]),
  .I1(ram16sdp_inst_876_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2341 (
  .O(mux_o_2341),
  .I0(ram16sdp_inst_884_dout[18]),
  .I1(ram16sdp_inst_892_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2342 (
  .O(mux_o_2342),
  .I0(ram16sdp_inst_900_dout[18]),
  .I1(ram16sdp_inst_908_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2343 (
  .O(mux_o_2343),
  .I0(ram16sdp_inst_916_dout[18]),
  .I1(ram16sdp_inst_924_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2344 (
  .O(mux_o_2344),
  .I0(ram16sdp_inst_932_dout[18]),
  .I1(ram16sdp_inst_940_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2345 (
  .O(mux_o_2345),
  .I0(ram16sdp_inst_948_dout[18]),
  .I1(ram16sdp_inst_956_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2346 (
  .O(mux_o_2346),
  .I0(ram16sdp_inst_964_dout[18]),
  .I1(ram16sdp_inst_972_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2347 (
  .O(mux_o_2347),
  .I0(ram16sdp_inst_980_dout[18]),
  .I1(ram16sdp_inst_988_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2348 (
  .O(mux_o_2348),
  .I0(ram16sdp_inst_996_dout[18]),
  .I1(ram16sdp_inst_1004_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2349 (
  .O(mux_o_2349),
  .I0(ram16sdp_inst_1012_dout[18]),
  .I1(ram16sdp_inst_1020_dout[18]),
  .S0(rad[4])
);
MUX2 mux_inst_2350 (
  .O(mux_o_2350),
  .I0(mux_o_2286),
  .I1(mux_o_2287),
  .S0(rad[5])
);
MUX2 mux_inst_2351 (
  .O(mux_o_2351),
  .I0(mux_o_2288),
  .I1(mux_o_2289),
  .S0(rad[5])
);
MUX2 mux_inst_2352 (
  .O(mux_o_2352),
  .I0(mux_o_2290),
  .I1(mux_o_2291),
  .S0(rad[5])
);
MUX2 mux_inst_2353 (
  .O(mux_o_2353),
  .I0(mux_o_2292),
  .I1(mux_o_2293),
  .S0(rad[5])
);
MUX2 mux_inst_2354 (
  .O(mux_o_2354),
  .I0(mux_o_2294),
  .I1(mux_o_2295),
  .S0(rad[5])
);
MUX2 mux_inst_2355 (
  .O(mux_o_2355),
  .I0(mux_o_2296),
  .I1(mux_o_2297),
  .S0(rad[5])
);
MUX2 mux_inst_2356 (
  .O(mux_o_2356),
  .I0(mux_o_2298),
  .I1(mux_o_2299),
  .S0(rad[5])
);
MUX2 mux_inst_2357 (
  .O(mux_o_2357),
  .I0(mux_o_2300),
  .I1(mux_o_2301),
  .S0(rad[5])
);
MUX2 mux_inst_2358 (
  .O(mux_o_2358),
  .I0(mux_o_2302),
  .I1(mux_o_2303),
  .S0(rad[5])
);
MUX2 mux_inst_2359 (
  .O(mux_o_2359),
  .I0(mux_o_2304),
  .I1(mux_o_2305),
  .S0(rad[5])
);
MUX2 mux_inst_2360 (
  .O(mux_o_2360),
  .I0(mux_o_2306),
  .I1(mux_o_2307),
  .S0(rad[5])
);
MUX2 mux_inst_2361 (
  .O(mux_o_2361),
  .I0(mux_o_2308),
  .I1(mux_o_2309),
  .S0(rad[5])
);
MUX2 mux_inst_2362 (
  .O(mux_o_2362),
  .I0(mux_o_2310),
  .I1(mux_o_2311),
  .S0(rad[5])
);
MUX2 mux_inst_2363 (
  .O(mux_o_2363),
  .I0(mux_o_2312),
  .I1(mux_o_2313),
  .S0(rad[5])
);
MUX2 mux_inst_2364 (
  .O(mux_o_2364),
  .I0(mux_o_2314),
  .I1(mux_o_2315),
  .S0(rad[5])
);
MUX2 mux_inst_2365 (
  .O(mux_o_2365),
  .I0(mux_o_2316),
  .I1(mux_o_2317),
  .S0(rad[5])
);
MUX2 mux_inst_2366 (
  .O(mux_o_2366),
  .I0(mux_o_2318),
  .I1(mux_o_2319),
  .S0(rad[5])
);
MUX2 mux_inst_2367 (
  .O(mux_o_2367),
  .I0(mux_o_2320),
  .I1(mux_o_2321),
  .S0(rad[5])
);
MUX2 mux_inst_2368 (
  .O(mux_o_2368),
  .I0(mux_o_2322),
  .I1(mux_o_2323),
  .S0(rad[5])
);
MUX2 mux_inst_2369 (
  .O(mux_o_2369),
  .I0(mux_o_2324),
  .I1(mux_o_2325),
  .S0(rad[5])
);
MUX2 mux_inst_2370 (
  .O(mux_o_2370),
  .I0(mux_o_2326),
  .I1(mux_o_2327),
  .S0(rad[5])
);
MUX2 mux_inst_2371 (
  .O(mux_o_2371),
  .I0(mux_o_2328),
  .I1(mux_o_2329),
  .S0(rad[5])
);
MUX2 mux_inst_2372 (
  .O(mux_o_2372),
  .I0(mux_o_2330),
  .I1(mux_o_2331),
  .S0(rad[5])
);
MUX2 mux_inst_2373 (
  .O(mux_o_2373),
  .I0(mux_o_2332),
  .I1(mux_o_2333),
  .S0(rad[5])
);
MUX2 mux_inst_2374 (
  .O(mux_o_2374),
  .I0(mux_o_2334),
  .I1(mux_o_2335),
  .S0(rad[5])
);
MUX2 mux_inst_2375 (
  .O(mux_o_2375),
  .I0(mux_o_2336),
  .I1(mux_o_2337),
  .S0(rad[5])
);
MUX2 mux_inst_2376 (
  .O(mux_o_2376),
  .I0(mux_o_2338),
  .I1(mux_o_2339),
  .S0(rad[5])
);
MUX2 mux_inst_2377 (
  .O(mux_o_2377),
  .I0(mux_o_2340),
  .I1(mux_o_2341),
  .S0(rad[5])
);
MUX2 mux_inst_2378 (
  .O(mux_o_2378),
  .I0(mux_o_2342),
  .I1(mux_o_2343),
  .S0(rad[5])
);
MUX2 mux_inst_2379 (
  .O(mux_o_2379),
  .I0(mux_o_2344),
  .I1(mux_o_2345),
  .S0(rad[5])
);
MUX2 mux_inst_2380 (
  .O(mux_o_2380),
  .I0(mux_o_2346),
  .I1(mux_o_2347),
  .S0(rad[5])
);
MUX2 mux_inst_2381 (
  .O(mux_o_2381),
  .I0(mux_o_2348),
  .I1(mux_o_2349),
  .S0(rad[5])
);
MUX2 mux_inst_2382 (
  .O(mux_o_2382),
  .I0(mux_o_2350),
  .I1(mux_o_2351),
  .S0(rad[6])
);
MUX2 mux_inst_2383 (
  .O(mux_o_2383),
  .I0(mux_o_2352),
  .I1(mux_o_2353),
  .S0(rad[6])
);
MUX2 mux_inst_2384 (
  .O(mux_o_2384),
  .I0(mux_o_2354),
  .I1(mux_o_2355),
  .S0(rad[6])
);
MUX2 mux_inst_2385 (
  .O(mux_o_2385),
  .I0(mux_o_2356),
  .I1(mux_o_2357),
  .S0(rad[6])
);
MUX2 mux_inst_2386 (
  .O(mux_o_2386),
  .I0(mux_o_2358),
  .I1(mux_o_2359),
  .S0(rad[6])
);
MUX2 mux_inst_2387 (
  .O(mux_o_2387),
  .I0(mux_o_2360),
  .I1(mux_o_2361),
  .S0(rad[6])
);
MUX2 mux_inst_2388 (
  .O(mux_o_2388),
  .I0(mux_o_2362),
  .I1(mux_o_2363),
  .S0(rad[6])
);
MUX2 mux_inst_2389 (
  .O(mux_o_2389),
  .I0(mux_o_2364),
  .I1(mux_o_2365),
  .S0(rad[6])
);
MUX2 mux_inst_2390 (
  .O(mux_o_2390),
  .I0(mux_o_2366),
  .I1(mux_o_2367),
  .S0(rad[6])
);
MUX2 mux_inst_2391 (
  .O(mux_o_2391),
  .I0(mux_o_2368),
  .I1(mux_o_2369),
  .S0(rad[6])
);
MUX2 mux_inst_2392 (
  .O(mux_o_2392),
  .I0(mux_o_2370),
  .I1(mux_o_2371),
  .S0(rad[6])
);
MUX2 mux_inst_2393 (
  .O(mux_o_2393),
  .I0(mux_o_2372),
  .I1(mux_o_2373),
  .S0(rad[6])
);
MUX2 mux_inst_2394 (
  .O(mux_o_2394),
  .I0(mux_o_2374),
  .I1(mux_o_2375),
  .S0(rad[6])
);
MUX2 mux_inst_2395 (
  .O(mux_o_2395),
  .I0(mux_o_2376),
  .I1(mux_o_2377),
  .S0(rad[6])
);
MUX2 mux_inst_2396 (
  .O(mux_o_2396),
  .I0(mux_o_2378),
  .I1(mux_o_2379),
  .S0(rad[6])
);
MUX2 mux_inst_2397 (
  .O(mux_o_2397),
  .I0(mux_o_2380),
  .I1(mux_o_2381),
  .S0(rad[6])
);
MUX2 mux_inst_2398 (
  .O(mux_o_2398),
  .I0(mux_o_2382),
  .I1(mux_o_2383),
  .S0(rad[7])
);
MUX2 mux_inst_2399 (
  .O(mux_o_2399),
  .I0(mux_o_2384),
  .I1(mux_o_2385),
  .S0(rad[7])
);
MUX2 mux_inst_2400 (
  .O(mux_o_2400),
  .I0(mux_o_2386),
  .I1(mux_o_2387),
  .S0(rad[7])
);
MUX2 mux_inst_2401 (
  .O(mux_o_2401),
  .I0(mux_o_2388),
  .I1(mux_o_2389),
  .S0(rad[7])
);
MUX2 mux_inst_2402 (
  .O(mux_o_2402),
  .I0(mux_o_2390),
  .I1(mux_o_2391),
  .S0(rad[7])
);
MUX2 mux_inst_2403 (
  .O(mux_o_2403),
  .I0(mux_o_2392),
  .I1(mux_o_2393),
  .S0(rad[7])
);
MUX2 mux_inst_2404 (
  .O(mux_o_2404),
  .I0(mux_o_2394),
  .I1(mux_o_2395),
  .S0(rad[7])
);
MUX2 mux_inst_2405 (
  .O(mux_o_2405),
  .I0(mux_o_2396),
  .I1(mux_o_2397),
  .S0(rad[7])
);
MUX2 mux_inst_2406 (
  .O(mux_o_2406),
  .I0(mux_o_2398),
  .I1(mux_o_2399),
  .S0(rad[8])
);
MUX2 mux_inst_2407 (
  .O(mux_o_2407),
  .I0(mux_o_2400),
  .I1(mux_o_2401),
  .S0(rad[8])
);
MUX2 mux_inst_2408 (
  .O(mux_o_2408),
  .I0(mux_o_2402),
  .I1(mux_o_2403),
  .S0(rad[8])
);
MUX2 mux_inst_2409 (
  .O(mux_o_2409),
  .I0(mux_o_2404),
  .I1(mux_o_2405),
  .S0(rad[8])
);
MUX2 mux_inst_2410 (
  .O(mux_o_2410),
  .I0(mux_o_2406),
  .I1(mux_o_2407),
  .S0(rad[9])
);
MUX2 mux_inst_2411 (
  .O(mux_o_2411),
  .I0(mux_o_2408),
  .I1(mux_o_2409),
  .S0(rad[9])
);
MUX2 mux_inst_2412 (
  .O(dout[18]),
  .I0(mux_o_2410),
  .I1(mux_o_2411),
  .S0(rad[10])
);
MUX2 mux_inst_2413 (
  .O(mux_o_2413),
  .I0(ram16sdp_inst_4_dout[19]),
  .I1(ram16sdp_inst_12_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2414 (
  .O(mux_o_2414),
  .I0(ram16sdp_inst_20_dout[19]),
  .I1(ram16sdp_inst_28_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2415 (
  .O(mux_o_2415),
  .I0(ram16sdp_inst_36_dout[19]),
  .I1(ram16sdp_inst_44_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2416 (
  .O(mux_o_2416),
  .I0(ram16sdp_inst_52_dout[19]),
  .I1(ram16sdp_inst_60_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2417 (
  .O(mux_o_2417),
  .I0(ram16sdp_inst_68_dout[19]),
  .I1(ram16sdp_inst_76_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2418 (
  .O(mux_o_2418),
  .I0(ram16sdp_inst_84_dout[19]),
  .I1(ram16sdp_inst_92_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2419 (
  .O(mux_o_2419),
  .I0(ram16sdp_inst_100_dout[19]),
  .I1(ram16sdp_inst_108_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2420 (
  .O(mux_o_2420),
  .I0(ram16sdp_inst_116_dout[19]),
  .I1(ram16sdp_inst_124_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2421 (
  .O(mux_o_2421),
  .I0(ram16sdp_inst_132_dout[19]),
  .I1(ram16sdp_inst_140_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2422 (
  .O(mux_o_2422),
  .I0(ram16sdp_inst_148_dout[19]),
  .I1(ram16sdp_inst_156_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2423 (
  .O(mux_o_2423),
  .I0(ram16sdp_inst_164_dout[19]),
  .I1(ram16sdp_inst_172_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2424 (
  .O(mux_o_2424),
  .I0(ram16sdp_inst_180_dout[19]),
  .I1(ram16sdp_inst_188_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2425 (
  .O(mux_o_2425),
  .I0(ram16sdp_inst_196_dout[19]),
  .I1(ram16sdp_inst_204_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2426 (
  .O(mux_o_2426),
  .I0(ram16sdp_inst_212_dout[19]),
  .I1(ram16sdp_inst_220_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2427 (
  .O(mux_o_2427),
  .I0(ram16sdp_inst_228_dout[19]),
  .I1(ram16sdp_inst_236_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2428 (
  .O(mux_o_2428),
  .I0(ram16sdp_inst_244_dout[19]),
  .I1(ram16sdp_inst_252_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2429 (
  .O(mux_o_2429),
  .I0(ram16sdp_inst_260_dout[19]),
  .I1(ram16sdp_inst_268_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2430 (
  .O(mux_o_2430),
  .I0(ram16sdp_inst_276_dout[19]),
  .I1(ram16sdp_inst_284_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2431 (
  .O(mux_o_2431),
  .I0(ram16sdp_inst_292_dout[19]),
  .I1(ram16sdp_inst_300_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2432 (
  .O(mux_o_2432),
  .I0(ram16sdp_inst_308_dout[19]),
  .I1(ram16sdp_inst_316_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2433 (
  .O(mux_o_2433),
  .I0(ram16sdp_inst_324_dout[19]),
  .I1(ram16sdp_inst_332_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2434 (
  .O(mux_o_2434),
  .I0(ram16sdp_inst_340_dout[19]),
  .I1(ram16sdp_inst_348_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2435 (
  .O(mux_o_2435),
  .I0(ram16sdp_inst_356_dout[19]),
  .I1(ram16sdp_inst_364_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2436 (
  .O(mux_o_2436),
  .I0(ram16sdp_inst_372_dout[19]),
  .I1(ram16sdp_inst_380_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2437 (
  .O(mux_o_2437),
  .I0(ram16sdp_inst_388_dout[19]),
  .I1(ram16sdp_inst_396_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2438 (
  .O(mux_o_2438),
  .I0(ram16sdp_inst_404_dout[19]),
  .I1(ram16sdp_inst_412_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2439 (
  .O(mux_o_2439),
  .I0(ram16sdp_inst_420_dout[19]),
  .I1(ram16sdp_inst_428_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2440 (
  .O(mux_o_2440),
  .I0(ram16sdp_inst_436_dout[19]),
  .I1(ram16sdp_inst_444_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2441 (
  .O(mux_o_2441),
  .I0(ram16sdp_inst_452_dout[19]),
  .I1(ram16sdp_inst_460_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2442 (
  .O(mux_o_2442),
  .I0(ram16sdp_inst_468_dout[19]),
  .I1(ram16sdp_inst_476_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2443 (
  .O(mux_o_2443),
  .I0(ram16sdp_inst_484_dout[19]),
  .I1(ram16sdp_inst_492_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2444 (
  .O(mux_o_2444),
  .I0(ram16sdp_inst_500_dout[19]),
  .I1(ram16sdp_inst_508_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2445 (
  .O(mux_o_2445),
  .I0(ram16sdp_inst_516_dout[19]),
  .I1(ram16sdp_inst_524_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2446 (
  .O(mux_o_2446),
  .I0(ram16sdp_inst_532_dout[19]),
  .I1(ram16sdp_inst_540_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2447 (
  .O(mux_o_2447),
  .I0(ram16sdp_inst_548_dout[19]),
  .I1(ram16sdp_inst_556_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2448 (
  .O(mux_o_2448),
  .I0(ram16sdp_inst_564_dout[19]),
  .I1(ram16sdp_inst_572_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2449 (
  .O(mux_o_2449),
  .I0(ram16sdp_inst_580_dout[19]),
  .I1(ram16sdp_inst_588_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2450 (
  .O(mux_o_2450),
  .I0(ram16sdp_inst_596_dout[19]),
  .I1(ram16sdp_inst_604_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2451 (
  .O(mux_o_2451),
  .I0(ram16sdp_inst_612_dout[19]),
  .I1(ram16sdp_inst_620_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2452 (
  .O(mux_o_2452),
  .I0(ram16sdp_inst_628_dout[19]),
  .I1(ram16sdp_inst_636_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2453 (
  .O(mux_o_2453),
  .I0(ram16sdp_inst_644_dout[19]),
  .I1(ram16sdp_inst_652_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2454 (
  .O(mux_o_2454),
  .I0(ram16sdp_inst_660_dout[19]),
  .I1(ram16sdp_inst_668_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2455 (
  .O(mux_o_2455),
  .I0(ram16sdp_inst_676_dout[19]),
  .I1(ram16sdp_inst_684_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2456 (
  .O(mux_o_2456),
  .I0(ram16sdp_inst_692_dout[19]),
  .I1(ram16sdp_inst_700_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2457 (
  .O(mux_o_2457),
  .I0(ram16sdp_inst_708_dout[19]),
  .I1(ram16sdp_inst_716_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2458 (
  .O(mux_o_2458),
  .I0(ram16sdp_inst_724_dout[19]),
  .I1(ram16sdp_inst_732_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2459 (
  .O(mux_o_2459),
  .I0(ram16sdp_inst_740_dout[19]),
  .I1(ram16sdp_inst_748_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2460 (
  .O(mux_o_2460),
  .I0(ram16sdp_inst_756_dout[19]),
  .I1(ram16sdp_inst_764_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2461 (
  .O(mux_o_2461),
  .I0(ram16sdp_inst_772_dout[19]),
  .I1(ram16sdp_inst_780_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2462 (
  .O(mux_o_2462),
  .I0(ram16sdp_inst_788_dout[19]),
  .I1(ram16sdp_inst_796_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2463 (
  .O(mux_o_2463),
  .I0(ram16sdp_inst_804_dout[19]),
  .I1(ram16sdp_inst_812_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2464 (
  .O(mux_o_2464),
  .I0(ram16sdp_inst_820_dout[19]),
  .I1(ram16sdp_inst_828_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2465 (
  .O(mux_o_2465),
  .I0(ram16sdp_inst_836_dout[19]),
  .I1(ram16sdp_inst_844_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2466 (
  .O(mux_o_2466),
  .I0(ram16sdp_inst_852_dout[19]),
  .I1(ram16sdp_inst_860_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2467 (
  .O(mux_o_2467),
  .I0(ram16sdp_inst_868_dout[19]),
  .I1(ram16sdp_inst_876_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2468 (
  .O(mux_o_2468),
  .I0(ram16sdp_inst_884_dout[19]),
  .I1(ram16sdp_inst_892_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2469 (
  .O(mux_o_2469),
  .I0(ram16sdp_inst_900_dout[19]),
  .I1(ram16sdp_inst_908_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2470 (
  .O(mux_o_2470),
  .I0(ram16sdp_inst_916_dout[19]),
  .I1(ram16sdp_inst_924_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2471 (
  .O(mux_o_2471),
  .I0(ram16sdp_inst_932_dout[19]),
  .I1(ram16sdp_inst_940_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2472 (
  .O(mux_o_2472),
  .I0(ram16sdp_inst_948_dout[19]),
  .I1(ram16sdp_inst_956_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2473 (
  .O(mux_o_2473),
  .I0(ram16sdp_inst_964_dout[19]),
  .I1(ram16sdp_inst_972_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2474 (
  .O(mux_o_2474),
  .I0(ram16sdp_inst_980_dout[19]),
  .I1(ram16sdp_inst_988_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2475 (
  .O(mux_o_2475),
  .I0(ram16sdp_inst_996_dout[19]),
  .I1(ram16sdp_inst_1004_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2476 (
  .O(mux_o_2476),
  .I0(ram16sdp_inst_1012_dout[19]),
  .I1(ram16sdp_inst_1020_dout[19]),
  .S0(rad[4])
);
MUX2 mux_inst_2477 (
  .O(mux_o_2477),
  .I0(mux_o_2413),
  .I1(mux_o_2414),
  .S0(rad[5])
);
MUX2 mux_inst_2478 (
  .O(mux_o_2478),
  .I0(mux_o_2415),
  .I1(mux_o_2416),
  .S0(rad[5])
);
MUX2 mux_inst_2479 (
  .O(mux_o_2479),
  .I0(mux_o_2417),
  .I1(mux_o_2418),
  .S0(rad[5])
);
MUX2 mux_inst_2480 (
  .O(mux_o_2480),
  .I0(mux_o_2419),
  .I1(mux_o_2420),
  .S0(rad[5])
);
MUX2 mux_inst_2481 (
  .O(mux_o_2481),
  .I0(mux_o_2421),
  .I1(mux_o_2422),
  .S0(rad[5])
);
MUX2 mux_inst_2482 (
  .O(mux_o_2482),
  .I0(mux_o_2423),
  .I1(mux_o_2424),
  .S0(rad[5])
);
MUX2 mux_inst_2483 (
  .O(mux_o_2483),
  .I0(mux_o_2425),
  .I1(mux_o_2426),
  .S0(rad[5])
);
MUX2 mux_inst_2484 (
  .O(mux_o_2484),
  .I0(mux_o_2427),
  .I1(mux_o_2428),
  .S0(rad[5])
);
MUX2 mux_inst_2485 (
  .O(mux_o_2485),
  .I0(mux_o_2429),
  .I1(mux_o_2430),
  .S0(rad[5])
);
MUX2 mux_inst_2486 (
  .O(mux_o_2486),
  .I0(mux_o_2431),
  .I1(mux_o_2432),
  .S0(rad[5])
);
MUX2 mux_inst_2487 (
  .O(mux_o_2487),
  .I0(mux_o_2433),
  .I1(mux_o_2434),
  .S0(rad[5])
);
MUX2 mux_inst_2488 (
  .O(mux_o_2488),
  .I0(mux_o_2435),
  .I1(mux_o_2436),
  .S0(rad[5])
);
MUX2 mux_inst_2489 (
  .O(mux_o_2489),
  .I0(mux_o_2437),
  .I1(mux_o_2438),
  .S0(rad[5])
);
MUX2 mux_inst_2490 (
  .O(mux_o_2490),
  .I0(mux_o_2439),
  .I1(mux_o_2440),
  .S0(rad[5])
);
MUX2 mux_inst_2491 (
  .O(mux_o_2491),
  .I0(mux_o_2441),
  .I1(mux_o_2442),
  .S0(rad[5])
);
MUX2 mux_inst_2492 (
  .O(mux_o_2492),
  .I0(mux_o_2443),
  .I1(mux_o_2444),
  .S0(rad[5])
);
MUX2 mux_inst_2493 (
  .O(mux_o_2493),
  .I0(mux_o_2445),
  .I1(mux_o_2446),
  .S0(rad[5])
);
MUX2 mux_inst_2494 (
  .O(mux_o_2494),
  .I0(mux_o_2447),
  .I1(mux_o_2448),
  .S0(rad[5])
);
MUX2 mux_inst_2495 (
  .O(mux_o_2495),
  .I0(mux_o_2449),
  .I1(mux_o_2450),
  .S0(rad[5])
);
MUX2 mux_inst_2496 (
  .O(mux_o_2496),
  .I0(mux_o_2451),
  .I1(mux_o_2452),
  .S0(rad[5])
);
MUX2 mux_inst_2497 (
  .O(mux_o_2497),
  .I0(mux_o_2453),
  .I1(mux_o_2454),
  .S0(rad[5])
);
MUX2 mux_inst_2498 (
  .O(mux_o_2498),
  .I0(mux_o_2455),
  .I1(mux_o_2456),
  .S0(rad[5])
);
MUX2 mux_inst_2499 (
  .O(mux_o_2499),
  .I0(mux_o_2457),
  .I1(mux_o_2458),
  .S0(rad[5])
);
MUX2 mux_inst_2500 (
  .O(mux_o_2500),
  .I0(mux_o_2459),
  .I1(mux_o_2460),
  .S0(rad[5])
);
MUX2 mux_inst_2501 (
  .O(mux_o_2501),
  .I0(mux_o_2461),
  .I1(mux_o_2462),
  .S0(rad[5])
);
MUX2 mux_inst_2502 (
  .O(mux_o_2502),
  .I0(mux_o_2463),
  .I1(mux_o_2464),
  .S0(rad[5])
);
MUX2 mux_inst_2503 (
  .O(mux_o_2503),
  .I0(mux_o_2465),
  .I1(mux_o_2466),
  .S0(rad[5])
);
MUX2 mux_inst_2504 (
  .O(mux_o_2504),
  .I0(mux_o_2467),
  .I1(mux_o_2468),
  .S0(rad[5])
);
MUX2 mux_inst_2505 (
  .O(mux_o_2505),
  .I0(mux_o_2469),
  .I1(mux_o_2470),
  .S0(rad[5])
);
MUX2 mux_inst_2506 (
  .O(mux_o_2506),
  .I0(mux_o_2471),
  .I1(mux_o_2472),
  .S0(rad[5])
);
MUX2 mux_inst_2507 (
  .O(mux_o_2507),
  .I0(mux_o_2473),
  .I1(mux_o_2474),
  .S0(rad[5])
);
MUX2 mux_inst_2508 (
  .O(mux_o_2508),
  .I0(mux_o_2475),
  .I1(mux_o_2476),
  .S0(rad[5])
);
MUX2 mux_inst_2509 (
  .O(mux_o_2509),
  .I0(mux_o_2477),
  .I1(mux_o_2478),
  .S0(rad[6])
);
MUX2 mux_inst_2510 (
  .O(mux_o_2510),
  .I0(mux_o_2479),
  .I1(mux_o_2480),
  .S0(rad[6])
);
MUX2 mux_inst_2511 (
  .O(mux_o_2511),
  .I0(mux_o_2481),
  .I1(mux_o_2482),
  .S0(rad[6])
);
MUX2 mux_inst_2512 (
  .O(mux_o_2512),
  .I0(mux_o_2483),
  .I1(mux_o_2484),
  .S0(rad[6])
);
MUX2 mux_inst_2513 (
  .O(mux_o_2513),
  .I0(mux_o_2485),
  .I1(mux_o_2486),
  .S0(rad[6])
);
MUX2 mux_inst_2514 (
  .O(mux_o_2514),
  .I0(mux_o_2487),
  .I1(mux_o_2488),
  .S0(rad[6])
);
MUX2 mux_inst_2515 (
  .O(mux_o_2515),
  .I0(mux_o_2489),
  .I1(mux_o_2490),
  .S0(rad[6])
);
MUX2 mux_inst_2516 (
  .O(mux_o_2516),
  .I0(mux_o_2491),
  .I1(mux_o_2492),
  .S0(rad[6])
);
MUX2 mux_inst_2517 (
  .O(mux_o_2517),
  .I0(mux_o_2493),
  .I1(mux_o_2494),
  .S0(rad[6])
);
MUX2 mux_inst_2518 (
  .O(mux_o_2518),
  .I0(mux_o_2495),
  .I1(mux_o_2496),
  .S0(rad[6])
);
MUX2 mux_inst_2519 (
  .O(mux_o_2519),
  .I0(mux_o_2497),
  .I1(mux_o_2498),
  .S0(rad[6])
);
MUX2 mux_inst_2520 (
  .O(mux_o_2520),
  .I0(mux_o_2499),
  .I1(mux_o_2500),
  .S0(rad[6])
);
MUX2 mux_inst_2521 (
  .O(mux_o_2521),
  .I0(mux_o_2501),
  .I1(mux_o_2502),
  .S0(rad[6])
);
MUX2 mux_inst_2522 (
  .O(mux_o_2522),
  .I0(mux_o_2503),
  .I1(mux_o_2504),
  .S0(rad[6])
);
MUX2 mux_inst_2523 (
  .O(mux_o_2523),
  .I0(mux_o_2505),
  .I1(mux_o_2506),
  .S0(rad[6])
);
MUX2 mux_inst_2524 (
  .O(mux_o_2524),
  .I0(mux_o_2507),
  .I1(mux_o_2508),
  .S0(rad[6])
);
MUX2 mux_inst_2525 (
  .O(mux_o_2525),
  .I0(mux_o_2509),
  .I1(mux_o_2510),
  .S0(rad[7])
);
MUX2 mux_inst_2526 (
  .O(mux_o_2526),
  .I0(mux_o_2511),
  .I1(mux_o_2512),
  .S0(rad[7])
);
MUX2 mux_inst_2527 (
  .O(mux_o_2527),
  .I0(mux_o_2513),
  .I1(mux_o_2514),
  .S0(rad[7])
);
MUX2 mux_inst_2528 (
  .O(mux_o_2528),
  .I0(mux_o_2515),
  .I1(mux_o_2516),
  .S0(rad[7])
);
MUX2 mux_inst_2529 (
  .O(mux_o_2529),
  .I0(mux_o_2517),
  .I1(mux_o_2518),
  .S0(rad[7])
);
MUX2 mux_inst_2530 (
  .O(mux_o_2530),
  .I0(mux_o_2519),
  .I1(mux_o_2520),
  .S0(rad[7])
);
MUX2 mux_inst_2531 (
  .O(mux_o_2531),
  .I0(mux_o_2521),
  .I1(mux_o_2522),
  .S0(rad[7])
);
MUX2 mux_inst_2532 (
  .O(mux_o_2532),
  .I0(mux_o_2523),
  .I1(mux_o_2524),
  .S0(rad[7])
);
MUX2 mux_inst_2533 (
  .O(mux_o_2533),
  .I0(mux_o_2525),
  .I1(mux_o_2526),
  .S0(rad[8])
);
MUX2 mux_inst_2534 (
  .O(mux_o_2534),
  .I0(mux_o_2527),
  .I1(mux_o_2528),
  .S0(rad[8])
);
MUX2 mux_inst_2535 (
  .O(mux_o_2535),
  .I0(mux_o_2529),
  .I1(mux_o_2530),
  .S0(rad[8])
);
MUX2 mux_inst_2536 (
  .O(mux_o_2536),
  .I0(mux_o_2531),
  .I1(mux_o_2532),
  .S0(rad[8])
);
MUX2 mux_inst_2537 (
  .O(mux_o_2537),
  .I0(mux_o_2533),
  .I1(mux_o_2534),
  .S0(rad[9])
);
MUX2 mux_inst_2538 (
  .O(mux_o_2538),
  .I0(mux_o_2535),
  .I1(mux_o_2536),
  .S0(rad[9])
);
MUX2 mux_inst_2539 (
  .O(dout[19]),
  .I0(mux_o_2537),
  .I1(mux_o_2538),
  .S0(rad[10])
);
MUX2 mux_inst_2540 (
  .O(mux_o_2540),
  .I0(ram16sdp_inst_5_dout[20]),
  .I1(ram16sdp_inst_13_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2541 (
  .O(mux_o_2541),
  .I0(ram16sdp_inst_21_dout[20]),
  .I1(ram16sdp_inst_29_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2542 (
  .O(mux_o_2542),
  .I0(ram16sdp_inst_37_dout[20]),
  .I1(ram16sdp_inst_45_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2543 (
  .O(mux_o_2543),
  .I0(ram16sdp_inst_53_dout[20]),
  .I1(ram16sdp_inst_61_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2544 (
  .O(mux_o_2544),
  .I0(ram16sdp_inst_69_dout[20]),
  .I1(ram16sdp_inst_77_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2545 (
  .O(mux_o_2545),
  .I0(ram16sdp_inst_85_dout[20]),
  .I1(ram16sdp_inst_93_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2546 (
  .O(mux_o_2546),
  .I0(ram16sdp_inst_101_dout[20]),
  .I1(ram16sdp_inst_109_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2547 (
  .O(mux_o_2547),
  .I0(ram16sdp_inst_117_dout[20]),
  .I1(ram16sdp_inst_125_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2548 (
  .O(mux_o_2548),
  .I0(ram16sdp_inst_133_dout[20]),
  .I1(ram16sdp_inst_141_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2549 (
  .O(mux_o_2549),
  .I0(ram16sdp_inst_149_dout[20]),
  .I1(ram16sdp_inst_157_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2550 (
  .O(mux_o_2550),
  .I0(ram16sdp_inst_165_dout[20]),
  .I1(ram16sdp_inst_173_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2551 (
  .O(mux_o_2551),
  .I0(ram16sdp_inst_181_dout[20]),
  .I1(ram16sdp_inst_189_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2552 (
  .O(mux_o_2552),
  .I0(ram16sdp_inst_197_dout[20]),
  .I1(ram16sdp_inst_205_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2553 (
  .O(mux_o_2553),
  .I0(ram16sdp_inst_213_dout[20]),
  .I1(ram16sdp_inst_221_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2554 (
  .O(mux_o_2554),
  .I0(ram16sdp_inst_229_dout[20]),
  .I1(ram16sdp_inst_237_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2555 (
  .O(mux_o_2555),
  .I0(ram16sdp_inst_245_dout[20]),
  .I1(ram16sdp_inst_253_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2556 (
  .O(mux_o_2556),
  .I0(ram16sdp_inst_261_dout[20]),
  .I1(ram16sdp_inst_269_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2557 (
  .O(mux_o_2557),
  .I0(ram16sdp_inst_277_dout[20]),
  .I1(ram16sdp_inst_285_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2558 (
  .O(mux_o_2558),
  .I0(ram16sdp_inst_293_dout[20]),
  .I1(ram16sdp_inst_301_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2559 (
  .O(mux_o_2559),
  .I0(ram16sdp_inst_309_dout[20]),
  .I1(ram16sdp_inst_317_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2560 (
  .O(mux_o_2560),
  .I0(ram16sdp_inst_325_dout[20]),
  .I1(ram16sdp_inst_333_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2561 (
  .O(mux_o_2561),
  .I0(ram16sdp_inst_341_dout[20]),
  .I1(ram16sdp_inst_349_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2562 (
  .O(mux_o_2562),
  .I0(ram16sdp_inst_357_dout[20]),
  .I1(ram16sdp_inst_365_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2563 (
  .O(mux_o_2563),
  .I0(ram16sdp_inst_373_dout[20]),
  .I1(ram16sdp_inst_381_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2564 (
  .O(mux_o_2564),
  .I0(ram16sdp_inst_389_dout[20]),
  .I1(ram16sdp_inst_397_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2565 (
  .O(mux_o_2565),
  .I0(ram16sdp_inst_405_dout[20]),
  .I1(ram16sdp_inst_413_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2566 (
  .O(mux_o_2566),
  .I0(ram16sdp_inst_421_dout[20]),
  .I1(ram16sdp_inst_429_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2567 (
  .O(mux_o_2567),
  .I0(ram16sdp_inst_437_dout[20]),
  .I1(ram16sdp_inst_445_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2568 (
  .O(mux_o_2568),
  .I0(ram16sdp_inst_453_dout[20]),
  .I1(ram16sdp_inst_461_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2569 (
  .O(mux_o_2569),
  .I0(ram16sdp_inst_469_dout[20]),
  .I1(ram16sdp_inst_477_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2570 (
  .O(mux_o_2570),
  .I0(ram16sdp_inst_485_dout[20]),
  .I1(ram16sdp_inst_493_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2571 (
  .O(mux_o_2571),
  .I0(ram16sdp_inst_501_dout[20]),
  .I1(ram16sdp_inst_509_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2572 (
  .O(mux_o_2572),
  .I0(ram16sdp_inst_517_dout[20]),
  .I1(ram16sdp_inst_525_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2573 (
  .O(mux_o_2573),
  .I0(ram16sdp_inst_533_dout[20]),
  .I1(ram16sdp_inst_541_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2574 (
  .O(mux_o_2574),
  .I0(ram16sdp_inst_549_dout[20]),
  .I1(ram16sdp_inst_557_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2575 (
  .O(mux_o_2575),
  .I0(ram16sdp_inst_565_dout[20]),
  .I1(ram16sdp_inst_573_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2576 (
  .O(mux_o_2576),
  .I0(ram16sdp_inst_581_dout[20]),
  .I1(ram16sdp_inst_589_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2577 (
  .O(mux_o_2577),
  .I0(ram16sdp_inst_597_dout[20]),
  .I1(ram16sdp_inst_605_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2578 (
  .O(mux_o_2578),
  .I0(ram16sdp_inst_613_dout[20]),
  .I1(ram16sdp_inst_621_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2579 (
  .O(mux_o_2579),
  .I0(ram16sdp_inst_629_dout[20]),
  .I1(ram16sdp_inst_637_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2580 (
  .O(mux_o_2580),
  .I0(ram16sdp_inst_645_dout[20]),
  .I1(ram16sdp_inst_653_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2581 (
  .O(mux_o_2581),
  .I0(ram16sdp_inst_661_dout[20]),
  .I1(ram16sdp_inst_669_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2582 (
  .O(mux_o_2582),
  .I0(ram16sdp_inst_677_dout[20]),
  .I1(ram16sdp_inst_685_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2583 (
  .O(mux_o_2583),
  .I0(ram16sdp_inst_693_dout[20]),
  .I1(ram16sdp_inst_701_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2584 (
  .O(mux_o_2584),
  .I0(ram16sdp_inst_709_dout[20]),
  .I1(ram16sdp_inst_717_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2585 (
  .O(mux_o_2585),
  .I0(ram16sdp_inst_725_dout[20]),
  .I1(ram16sdp_inst_733_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2586 (
  .O(mux_o_2586),
  .I0(ram16sdp_inst_741_dout[20]),
  .I1(ram16sdp_inst_749_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2587 (
  .O(mux_o_2587),
  .I0(ram16sdp_inst_757_dout[20]),
  .I1(ram16sdp_inst_765_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2588 (
  .O(mux_o_2588),
  .I0(ram16sdp_inst_773_dout[20]),
  .I1(ram16sdp_inst_781_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2589 (
  .O(mux_o_2589),
  .I0(ram16sdp_inst_789_dout[20]),
  .I1(ram16sdp_inst_797_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2590 (
  .O(mux_o_2590),
  .I0(ram16sdp_inst_805_dout[20]),
  .I1(ram16sdp_inst_813_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2591 (
  .O(mux_o_2591),
  .I0(ram16sdp_inst_821_dout[20]),
  .I1(ram16sdp_inst_829_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2592 (
  .O(mux_o_2592),
  .I0(ram16sdp_inst_837_dout[20]),
  .I1(ram16sdp_inst_845_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2593 (
  .O(mux_o_2593),
  .I0(ram16sdp_inst_853_dout[20]),
  .I1(ram16sdp_inst_861_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2594 (
  .O(mux_o_2594),
  .I0(ram16sdp_inst_869_dout[20]),
  .I1(ram16sdp_inst_877_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2595 (
  .O(mux_o_2595),
  .I0(ram16sdp_inst_885_dout[20]),
  .I1(ram16sdp_inst_893_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2596 (
  .O(mux_o_2596),
  .I0(ram16sdp_inst_901_dout[20]),
  .I1(ram16sdp_inst_909_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2597 (
  .O(mux_o_2597),
  .I0(ram16sdp_inst_917_dout[20]),
  .I1(ram16sdp_inst_925_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2598 (
  .O(mux_o_2598),
  .I0(ram16sdp_inst_933_dout[20]),
  .I1(ram16sdp_inst_941_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2599 (
  .O(mux_o_2599),
  .I0(ram16sdp_inst_949_dout[20]),
  .I1(ram16sdp_inst_957_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2600 (
  .O(mux_o_2600),
  .I0(ram16sdp_inst_965_dout[20]),
  .I1(ram16sdp_inst_973_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2601 (
  .O(mux_o_2601),
  .I0(ram16sdp_inst_981_dout[20]),
  .I1(ram16sdp_inst_989_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2602 (
  .O(mux_o_2602),
  .I0(ram16sdp_inst_997_dout[20]),
  .I1(ram16sdp_inst_1005_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2603 (
  .O(mux_o_2603),
  .I0(ram16sdp_inst_1013_dout[20]),
  .I1(ram16sdp_inst_1021_dout[20]),
  .S0(rad[4])
);
MUX2 mux_inst_2604 (
  .O(mux_o_2604),
  .I0(mux_o_2540),
  .I1(mux_o_2541),
  .S0(rad[5])
);
MUX2 mux_inst_2605 (
  .O(mux_o_2605),
  .I0(mux_o_2542),
  .I1(mux_o_2543),
  .S0(rad[5])
);
MUX2 mux_inst_2606 (
  .O(mux_o_2606),
  .I0(mux_o_2544),
  .I1(mux_o_2545),
  .S0(rad[5])
);
MUX2 mux_inst_2607 (
  .O(mux_o_2607),
  .I0(mux_o_2546),
  .I1(mux_o_2547),
  .S0(rad[5])
);
MUX2 mux_inst_2608 (
  .O(mux_o_2608),
  .I0(mux_o_2548),
  .I1(mux_o_2549),
  .S0(rad[5])
);
MUX2 mux_inst_2609 (
  .O(mux_o_2609),
  .I0(mux_o_2550),
  .I1(mux_o_2551),
  .S0(rad[5])
);
MUX2 mux_inst_2610 (
  .O(mux_o_2610),
  .I0(mux_o_2552),
  .I1(mux_o_2553),
  .S0(rad[5])
);
MUX2 mux_inst_2611 (
  .O(mux_o_2611),
  .I0(mux_o_2554),
  .I1(mux_o_2555),
  .S0(rad[5])
);
MUX2 mux_inst_2612 (
  .O(mux_o_2612),
  .I0(mux_o_2556),
  .I1(mux_o_2557),
  .S0(rad[5])
);
MUX2 mux_inst_2613 (
  .O(mux_o_2613),
  .I0(mux_o_2558),
  .I1(mux_o_2559),
  .S0(rad[5])
);
MUX2 mux_inst_2614 (
  .O(mux_o_2614),
  .I0(mux_o_2560),
  .I1(mux_o_2561),
  .S0(rad[5])
);
MUX2 mux_inst_2615 (
  .O(mux_o_2615),
  .I0(mux_o_2562),
  .I1(mux_o_2563),
  .S0(rad[5])
);
MUX2 mux_inst_2616 (
  .O(mux_o_2616),
  .I0(mux_o_2564),
  .I1(mux_o_2565),
  .S0(rad[5])
);
MUX2 mux_inst_2617 (
  .O(mux_o_2617),
  .I0(mux_o_2566),
  .I1(mux_o_2567),
  .S0(rad[5])
);
MUX2 mux_inst_2618 (
  .O(mux_o_2618),
  .I0(mux_o_2568),
  .I1(mux_o_2569),
  .S0(rad[5])
);
MUX2 mux_inst_2619 (
  .O(mux_o_2619),
  .I0(mux_o_2570),
  .I1(mux_o_2571),
  .S0(rad[5])
);
MUX2 mux_inst_2620 (
  .O(mux_o_2620),
  .I0(mux_o_2572),
  .I1(mux_o_2573),
  .S0(rad[5])
);
MUX2 mux_inst_2621 (
  .O(mux_o_2621),
  .I0(mux_o_2574),
  .I1(mux_o_2575),
  .S0(rad[5])
);
MUX2 mux_inst_2622 (
  .O(mux_o_2622),
  .I0(mux_o_2576),
  .I1(mux_o_2577),
  .S0(rad[5])
);
MUX2 mux_inst_2623 (
  .O(mux_o_2623),
  .I0(mux_o_2578),
  .I1(mux_o_2579),
  .S0(rad[5])
);
MUX2 mux_inst_2624 (
  .O(mux_o_2624),
  .I0(mux_o_2580),
  .I1(mux_o_2581),
  .S0(rad[5])
);
MUX2 mux_inst_2625 (
  .O(mux_o_2625),
  .I0(mux_o_2582),
  .I1(mux_o_2583),
  .S0(rad[5])
);
MUX2 mux_inst_2626 (
  .O(mux_o_2626),
  .I0(mux_o_2584),
  .I1(mux_o_2585),
  .S0(rad[5])
);
MUX2 mux_inst_2627 (
  .O(mux_o_2627),
  .I0(mux_o_2586),
  .I1(mux_o_2587),
  .S0(rad[5])
);
MUX2 mux_inst_2628 (
  .O(mux_o_2628),
  .I0(mux_o_2588),
  .I1(mux_o_2589),
  .S0(rad[5])
);
MUX2 mux_inst_2629 (
  .O(mux_o_2629),
  .I0(mux_o_2590),
  .I1(mux_o_2591),
  .S0(rad[5])
);
MUX2 mux_inst_2630 (
  .O(mux_o_2630),
  .I0(mux_o_2592),
  .I1(mux_o_2593),
  .S0(rad[5])
);
MUX2 mux_inst_2631 (
  .O(mux_o_2631),
  .I0(mux_o_2594),
  .I1(mux_o_2595),
  .S0(rad[5])
);
MUX2 mux_inst_2632 (
  .O(mux_o_2632),
  .I0(mux_o_2596),
  .I1(mux_o_2597),
  .S0(rad[5])
);
MUX2 mux_inst_2633 (
  .O(mux_o_2633),
  .I0(mux_o_2598),
  .I1(mux_o_2599),
  .S0(rad[5])
);
MUX2 mux_inst_2634 (
  .O(mux_o_2634),
  .I0(mux_o_2600),
  .I1(mux_o_2601),
  .S0(rad[5])
);
MUX2 mux_inst_2635 (
  .O(mux_o_2635),
  .I0(mux_o_2602),
  .I1(mux_o_2603),
  .S0(rad[5])
);
MUX2 mux_inst_2636 (
  .O(mux_o_2636),
  .I0(mux_o_2604),
  .I1(mux_o_2605),
  .S0(rad[6])
);
MUX2 mux_inst_2637 (
  .O(mux_o_2637),
  .I0(mux_o_2606),
  .I1(mux_o_2607),
  .S0(rad[6])
);
MUX2 mux_inst_2638 (
  .O(mux_o_2638),
  .I0(mux_o_2608),
  .I1(mux_o_2609),
  .S0(rad[6])
);
MUX2 mux_inst_2639 (
  .O(mux_o_2639),
  .I0(mux_o_2610),
  .I1(mux_o_2611),
  .S0(rad[6])
);
MUX2 mux_inst_2640 (
  .O(mux_o_2640),
  .I0(mux_o_2612),
  .I1(mux_o_2613),
  .S0(rad[6])
);
MUX2 mux_inst_2641 (
  .O(mux_o_2641),
  .I0(mux_o_2614),
  .I1(mux_o_2615),
  .S0(rad[6])
);
MUX2 mux_inst_2642 (
  .O(mux_o_2642),
  .I0(mux_o_2616),
  .I1(mux_o_2617),
  .S0(rad[6])
);
MUX2 mux_inst_2643 (
  .O(mux_o_2643),
  .I0(mux_o_2618),
  .I1(mux_o_2619),
  .S0(rad[6])
);
MUX2 mux_inst_2644 (
  .O(mux_o_2644),
  .I0(mux_o_2620),
  .I1(mux_o_2621),
  .S0(rad[6])
);
MUX2 mux_inst_2645 (
  .O(mux_o_2645),
  .I0(mux_o_2622),
  .I1(mux_o_2623),
  .S0(rad[6])
);
MUX2 mux_inst_2646 (
  .O(mux_o_2646),
  .I0(mux_o_2624),
  .I1(mux_o_2625),
  .S0(rad[6])
);
MUX2 mux_inst_2647 (
  .O(mux_o_2647),
  .I0(mux_o_2626),
  .I1(mux_o_2627),
  .S0(rad[6])
);
MUX2 mux_inst_2648 (
  .O(mux_o_2648),
  .I0(mux_o_2628),
  .I1(mux_o_2629),
  .S0(rad[6])
);
MUX2 mux_inst_2649 (
  .O(mux_o_2649),
  .I0(mux_o_2630),
  .I1(mux_o_2631),
  .S0(rad[6])
);
MUX2 mux_inst_2650 (
  .O(mux_o_2650),
  .I0(mux_o_2632),
  .I1(mux_o_2633),
  .S0(rad[6])
);
MUX2 mux_inst_2651 (
  .O(mux_o_2651),
  .I0(mux_o_2634),
  .I1(mux_o_2635),
  .S0(rad[6])
);
MUX2 mux_inst_2652 (
  .O(mux_o_2652),
  .I0(mux_o_2636),
  .I1(mux_o_2637),
  .S0(rad[7])
);
MUX2 mux_inst_2653 (
  .O(mux_o_2653),
  .I0(mux_o_2638),
  .I1(mux_o_2639),
  .S0(rad[7])
);
MUX2 mux_inst_2654 (
  .O(mux_o_2654),
  .I0(mux_o_2640),
  .I1(mux_o_2641),
  .S0(rad[7])
);
MUX2 mux_inst_2655 (
  .O(mux_o_2655),
  .I0(mux_o_2642),
  .I1(mux_o_2643),
  .S0(rad[7])
);
MUX2 mux_inst_2656 (
  .O(mux_o_2656),
  .I0(mux_o_2644),
  .I1(mux_o_2645),
  .S0(rad[7])
);
MUX2 mux_inst_2657 (
  .O(mux_o_2657),
  .I0(mux_o_2646),
  .I1(mux_o_2647),
  .S0(rad[7])
);
MUX2 mux_inst_2658 (
  .O(mux_o_2658),
  .I0(mux_o_2648),
  .I1(mux_o_2649),
  .S0(rad[7])
);
MUX2 mux_inst_2659 (
  .O(mux_o_2659),
  .I0(mux_o_2650),
  .I1(mux_o_2651),
  .S0(rad[7])
);
MUX2 mux_inst_2660 (
  .O(mux_o_2660),
  .I0(mux_o_2652),
  .I1(mux_o_2653),
  .S0(rad[8])
);
MUX2 mux_inst_2661 (
  .O(mux_o_2661),
  .I0(mux_o_2654),
  .I1(mux_o_2655),
  .S0(rad[8])
);
MUX2 mux_inst_2662 (
  .O(mux_o_2662),
  .I0(mux_o_2656),
  .I1(mux_o_2657),
  .S0(rad[8])
);
MUX2 mux_inst_2663 (
  .O(mux_o_2663),
  .I0(mux_o_2658),
  .I1(mux_o_2659),
  .S0(rad[8])
);
MUX2 mux_inst_2664 (
  .O(mux_o_2664),
  .I0(mux_o_2660),
  .I1(mux_o_2661),
  .S0(rad[9])
);
MUX2 mux_inst_2665 (
  .O(mux_o_2665),
  .I0(mux_o_2662),
  .I1(mux_o_2663),
  .S0(rad[9])
);
MUX2 mux_inst_2666 (
  .O(dout[20]),
  .I0(mux_o_2664),
  .I1(mux_o_2665),
  .S0(rad[10])
);
MUX2 mux_inst_2667 (
  .O(mux_o_2667),
  .I0(ram16sdp_inst_5_dout[21]),
  .I1(ram16sdp_inst_13_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2668 (
  .O(mux_o_2668),
  .I0(ram16sdp_inst_21_dout[21]),
  .I1(ram16sdp_inst_29_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2669 (
  .O(mux_o_2669),
  .I0(ram16sdp_inst_37_dout[21]),
  .I1(ram16sdp_inst_45_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2670 (
  .O(mux_o_2670),
  .I0(ram16sdp_inst_53_dout[21]),
  .I1(ram16sdp_inst_61_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2671 (
  .O(mux_o_2671),
  .I0(ram16sdp_inst_69_dout[21]),
  .I1(ram16sdp_inst_77_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2672 (
  .O(mux_o_2672),
  .I0(ram16sdp_inst_85_dout[21]),
  .I1(ram16sdp_inst_93_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2673 (
  .O(mux_o_2673),
  .I0(ram16sdp_inst_101_dout[21]),
  .I1(ram16sdp_inst_109_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2674 (
  .O(mux_o_2674),
  .I0(ram16sdp_inst_117_dout[21]),
  .I1(ram16sdp_inst_125_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2675 (
  .O(mux_o_2675),
  .I0(ram16sdp_inst_133_dout[21]),
  .I1(ram16sdp_inst_141_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2676 (
  .O(mux_o_2676),
  .I0(ram16sdp_inst_149_dout[21]),
  .I1(ram16sdp_inst_157_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2677 (
  .O(mux_o_2677),
  .I0(ram16sdp_inst_165_dout[21]),
  .I1(ram16sdp_inst_173_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2678 (
  .O(mux_o_2678),
  .I0(ram16sdp_inst_181_dout[21]),
  .I1(ram16sdp_inst_189_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2679 (
  .O(mux_o_2679),
  .I0(ram16sdp_inst_197_dout[21]),
  .I1(ram16sdp_inst_205_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2680 (
  .O(mux_o_2680),
  .I0(ram16sdp_inst_213_dout[21]),
  .I1(ram16sdp_inst_221_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2681 (
  .O(mux_o_2681),
  .I0(ram16sdp_inst_229_dout[21]),
  .I1(ram16sdp_inst_237_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2682 (
  .O(mux_o_2682),
  .I0(ram16sdp_inst_245_dout[21]),
  .I1(ram16sdp_inst_253_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2683 (
  .O(mux_o_2683),
  .I0(ram16sdp_inst_261_dout[21]),
  .I1(ram16sdp_inst_269_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2684 (
  .O(mux_o_2684),
  .I0(ram16sdp_inst_277_dout[21]),
  .I1(ram16sdp_inst_285_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2685 (
  .O(mux_o_2685),
  .I0(ram16sdp_inst_293_dout[21]),
  .I1(ram16sdp_inst_301_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2686 (
  .O(mux_o_2686),
  .I0(ram16sdp_inst_309_dout[21]),
  .I1(ram16sdp_inst_317_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2687 (
  .O(mux_o_2687),
  .I0(ram16sdp_inst_325_dout[21]),
  .I1(ram16sdp_inst_333_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2688 (
  .O(mux_o_2688),
  .I0(ram16sdp_inst_341_dout[21]),
  .I1(ram16sdp_inst_349_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2689 (
  .O(mux_o_2689),
  .I0(ram16sdp_inst_357_dout[21]),
  .I1(ram16sdp_inst_365_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2690 (
  .O(mux_o_2690),
  .I0(ram16sdp_inst_373_dout[21]),
  .I1(ram16sdp_inst_381_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2691 (
  .O(mux_o_2691),
  .I0(ram16sdp_inst_389_dout[21]),
  .I1(ram16sdp_inst_397_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2692 (
  .O(mux_o_2692),
  .I0(ram16sdp_inst_405_dout[21]),
  .I1(ram16sdp_inst_413_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2693 (
  .O(mux_o_2693),
  .I0(ram16sdp_inst_421_dout[21]),
  .I1(ram16sdp_inst_429_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2694 (
  .O(mux_o_2694),
  .I0(ram16sdp_inst_437_dout[21]),
  .I1(ram16sdp_inst_445_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2695 (
  .O(mux_o_2695),
  .I0(ram16sdp_inst_453_dout[21]),
  .I1(ram16sdp_inst_461_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2696 (
  .O(mux_o_2696),
  .I0(ram16sdp_inst_469_dout[21]),
  .I1(ram16sdp_inst_477_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2697 (
  .O(mux_o_2697),
  .I0(ram16sdp_inst_485_dout[21]),
  .I1(ram16sdp_inst_493_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2698 (
  .O(mux_o_2698),
  .I0(ram16sdp_inst_501_dout[21]),
  .I1(ram16sdp_inst_509_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2699 (
  .O(mux_o_2699),
  .I0(ram16sdp_inst_517_dout[21]),
  .I1(ram16sdp_inst_525_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2700 (
  .O(mux_o_2700),
  .I0(ram16sdp_inst_533_dout[21]),
  .I1(ram16sdp_inst_541_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2701 (
  .O(mux_o_2701),
  .I0(ram16sdp_inst_549_dout[21]),
  .I1(ram16sdp_inst_557_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2702 (
  .O(mux_o_2702),
  .I0(ram16sdp_inst_565_dout[21]),
  .I1(ram16sdp_inst_573_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2703 (
  .O(mux_o_2703),
  .I0(ram16sdp_inst_581_dout[21]),
  .I1(ram16sdp_inst_589_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2704 (
  .O(mux_o_2704),
  .I0(ram16sdp_inst_597_dout[21]),
  .I1(ram16sdp_inst_605_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2705 (
  .O(mux_o_2705),
  .I0(ram16sdp_inst_613_dout[21]),
  .I1(ram16sdp_inst_621_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2706 (
  .O(mux_o_2706),
  .I0(ram16sdp_inst_629_dout[21]),
  .I1(ram16sdp_inst_637_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2707 (
  .O(mux_o_2707),
  .I0(ram16sdp_inst_645_dout[21]),
  .I1(ram16sdp_inst_653_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2708 (
  .O(mux_o_2708),
  .I0(ram16sdp_inst_661_dout[21]),
  .I1(ram16sdp_inst_669_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2709 (
  .O(mux_o_2709),
  .I0(ram16sdp_inst_677_dout[21]),
  .I1(ram16sdp_inst_685_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2710 (
  .O(mux_o_2710),
  .I0(ram16sdp_inst_693_dout[21]),
  .I1(ram16sdp_inst_701_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2711 (
  .O(mux_o_2711),
  .I0(ram16sdp_inst_709_dout[21]),
  .I1(ram16sdp_inst_717_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2712 (
  .O(mux_o_2712),
  .I0(ram16sdp_inst_725_dout[21]),
  .I1(ram16sdp_inst_733_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2713 (
  .O(mux_o_2713),
  .I0(ram16sdp_inst_741_dout[21]),
  .I1(ram16sdp_inst_749_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2714 (
  .O(mux_o_2714),
  .I0(ram16sdp_inst_757_dout[21]),
  .I1(ram16sdp_inst_765_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2715 (
  .O(mux_o_2715),
  .I0(ram16sdp_inst_773_dout[21]),
  .I1(ram16sdp_inst_781_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2716 (
  .O(mux_o_2716),
  .I0(ram16sdp_inst_789_dout[21]),
  .I1(ram16sdp_inst_797_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2717 (
  .O(mux_o_2717),
  .I0(ram16sdp_inst_805_dout[21]),
  .I1(ram16sdp_inst_813_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2718 (
  .O(mux_o_2718),
  .I0(ram16sdp_inst_821_dout[21]),
  .I1(ram16sdp_inst_829_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2719 (
  .O(mux_o_2719),
  .I0(ram16sdp_inst_837_dout[21]),
  .I1(ram16sdp_inst_845_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2720 (
  .O(mux_o_2720),
  .I0(ram16sdp_inst_853_dout[21]),
  .I1(ram16sdp_inst_861_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2721 (
  .O(mux_o_2721),
  .I0(ram16sdp_inst_869_dout[21]),
  .I1(ram16sdp_inst_877_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2722 (
  .O(mux_o_2722),
  .I0(ram16sdp_inst_885_dout[21]),
  .I1(ram16sdp_inst_893_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2723 (
  .O(mux_o_2723),
  .I0(ram16sdp_inst_901_dout[21]),
  .I1(ram16sdp_inst_909_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2724 (
  .O(mux_o_2724),
  .I0(ram16sdp_inst_917_dout[21]),
  .I1(ram16sdp_inst_925_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2725 (
  .O(mux_o_2725),
  .I0(ram16sdp_inst_933_dout[21]),
  .I1(ram16sdp_inst_941_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2726 (
  .O(mux_o_2726),
  .I0(ram16sdp_inst_949_dout[21]),
  .I1(ram16sdp_inst_957_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2727 (
  .O(mux_o_2727),
  .I0(ram16sdp_inst_965_dout[21]),
  .I1(ram16sdp_inst_973_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2728 (
  .O(mux_o_2728),
  .I0(ram16sdp_inst_981_dout[21]),
  .I1(ram16sdp_inst_989_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2729 (
  .O(mux_o_2729),
  .I0(ram16sdp_inst_997_dout[21]),
  .I1(ram16sdp_inst_1005_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2730 (
  .O(mux_o_2730),
  .I0(ram16sdp_inst_1013_dout[21]),
  .I1(ram16sdp_inst_1021_dout[21]),
  .S0(rad[4])
);
MUX2 mux_inst_2731 (
  .O(mux_o_2731),
  .I0(mux_o_2667),
  .I1(mux_o_2668),
  .S0(rad[5])
);
MUX2 mux_inst_2732 (
  .O(mux_o_2732),
  .I0(mux_o_2669),
  .I1(mux_o_2670),
  .S0(rad[5])
);
MUX2 mux_inst_2733 (
  .O(mux_o_2733),
  .I0(mux_o_2671),
  .I1(mux_o_2672),
  .S0(rad[5])
);
MUX2 mux_inst_2734 (
  .O(mux_o_2734),
  .I0(mux_o_2673),
  .I1(mux_o_2674),
  .S0(rad[5])
);
MUX2 mux_inst_2735 (
  .O(mux_o_2735),
  .I0(mux_o_2675),
  .I1(mux_o_2676),
  .S0(rad[5])
);
MUX2 mux_inst_2736 (
  .O(mux_o_2736),
  .I0(mux_o_2677),
  .I1(mux_o_2678),
  .S0(rad[5])
);
MUX2 mux_inst_2737 (
  .O(mux_o_2737),
  .I0(mux_o_2679),
  .I1(mux_o_2680),
  .S0(rad[5])
);
MUX2 mux_inst_2738 (
  .O(mux_o_2738),
  .I0(mux_o_2681),
  .I1(mux_o_2682),
  .S0(rad[5])
);
MUX2 mux_inst_2739 (
  .O(mux_o_2739),
  .I0(mux_o_2683),
  .I1(mux_o_2684),
  .S0(rad[5])
);
MUX2 mux_inst_2740 (
  .O(mux_o_2740),
  .I0(mux_o_2685),
  .I1(mux_o_2686),
  .S0(rad[5])
);
MUX2 mux_inst_2741 (
  .O(mux_o_2741),
  .I0(mux_o_2687),
  .I1(mux_o_2688),
  .S0(rad[5])
);
MUX2 mux_inst_2742 (
  .O(mux_o_2742),
  .I0(mux_o_2689),
  .I1(mux_o_2690),
  .S0(rad[5])
);
MUX2 mux_inst_2743 (
  .O(mux_o_2743),
  .I0(mux_o_2691),
  .I1(mux_o_2692),
  .S0(rad[5])
);
MUX2 mux_inst_2744 (
  .O(mux_o_2744),
  .I0(mux_o_2693),
  .I1(mux_o_2694),
  .S0(rad[5])
);
MUX2 mux_inst_2745 (
  .O(mux_o_2745),
  .I0(mux_o_2695),
  .I1(mux_o_2696),
  .S0(rad[5])
);
MUX2 mux_inst_2746 (
  .O(mux_o_2746),
  .I0(mux_o_2697),
  .I1(mux_o_2698),
  .S0(rad[5])
);
MUX2 mux_inst_2747 (
  .O(mux_o_2747),
  .I0(mux_o_2699),
  .I1(mux_o_2700),
  .S0(rad[5])
);
MUX2 mux_inst_2748 (
  .O(mux_o_2748),
  .I0(mux_o_2701),
  .I1(mux_o_2702),
  .S0(rad[5])
);
MUX2 mux_inst_2749 (
  .O(mux_o_2749),
  .I0(mux_o_2703),
  .I1(mux_o_2704),
  .S0(rad[5])
);
MUX2 mux_inst_2750 (
  .O(mux_o_2750),
  .I0(mux_o_2705),
  .I1(mux_o_2706),
  .S0(rad[5])
);
MUX2 mux_inst_2751 (
  .O(mux_o_2751),
  .I0(mux_o_2707),
  .I1(mux_o_2708),
  .S0(rad[5])
);
MUX2 mux_inst_2752 (
  .O(mux_o_2752),
  .I0(mux_o_2709),
  .I1(mux_o_2710),
  .S0(rad[5])
);
MUX2 mux_inst_2753 (
  .O(mux_o_2753),
  .I0(mux_o_2711),
  .I1(mux_o_2712),
  .S0(rad[5])
);
MUX2 mux_inst_2754 (
  .O(mux_o_2754),
  .I0(mux_o_2713),
  .I1(mux_o_2714),
  .S0(rad[5])
);
MUX2 mux_inst_2755 (
  .O(mux_o_2755),
  .I0(mux_o_2715),
  .I1(mux_o_2716),
  .S0(rad[5])
);
MUX2 mux_inst_2756 (
  .O(mux_o_2756),
  .I0(mux_o_2717),
  .I1(mux_o_2718),
  .S0(rad[5])
);
MUX2 mux_inst_2757 (
  .O(mux_o_2757),
  .I0(mux_o_2719),
  .I1(mux_o_2720),
  .S0(rad[5])
);
MUX2 mux_inst_2758 (
  .O(mux_o_2758),
  .I0(mux_o_2721),
  .I1(mux_o_2722),
  .S0(rad[5])
);
MUX2 mux_inst_2759 (
  .O(mux_o_2759),
  .I0(mux_o_2723),
  .I1(mux_o_2724),
  .S0(rad[5])
);
MUX2 mux_inst_2760 (
  .O(mux_o_2760),
  .I0(mux_o_2725),
  .I1(mux_o_2726),
  .S0(rad[5])
);
MUX2 mux_inst_2761 (
  .O(mux_o_2761),
  .I0(mux_o_2727),
  .I1(mux_o_2728),
  .S0(rad[5])
);
MUX2 mux_inst_2762 (
  .O(mux_o_2762),
  .I0(mux_o_2729),
  .I1(mux_o_2730),
  .S0(rad[5])
);
MUX2 mux_inst_2763 (
  .O(mux_o_2763),
  .I0(mux_o_2731),
  .I1(mux_o_2732),
  .S0(rad[6])
);
MUX2 mux_inst_2764 (
  .O(mux_o_2764),
  .I0(mux_o_2733),
  .I1(mux_o_2734),
  .S0(rad[6])
);
MUX2 mux_inst_2765 (
  .O(mux_o_2765),
  .I0(mux_o_2735),
  .I1(mux_o_2736),
  .S0(rad[6])
);
MUX2 mux_inst_2766 (
  .O(mux_o_2766),
  .I0(mux_o_2737),
  .I1(mux_o_2738),
  .S0(rad[6])
);
MUX2 mux_inst_2767 (
  .O(mux_o_2767),
  .I0(mux_o_2739),
  .I1(mux_o_2740),
  .S0(rad[6])
);
MUX2 mux_inst_2768 (
  .O(mux_o_2768),
  .I0(mux_o_2741),
  .I1(mux_o_2742),
  .S0(rad[6])
);
MUX2 mux_inst_2769 (
  .O(mux_o_2769),
  .I0(mux_o_2743),
  .I1(mux_o_2744),
  .S0(rad[6])
);
MUX2 mux_inst_2770 (
  .O(mux_o_2770),
  .I0(mux_o_2745),
  .I1(mux_o_2746),
  .S0(rad[6])
);
MUX2 mux_inst_2771 (
  .O(mux_o_2771),
  .I0(mux_o_2747),
  .I1(mux_o_2748),
  .S0(rad[6])
);
MUX2 mux_inst_2772 (
  .O(mux_o_2772),
  .I0(mux_o_2749),
  .I1(mux_o_2750),
  .S0(rad[6])
);
MUX2 mux_inst_2773 (
  .O(mux_o_2773),
  .I0(mux_o_2751),
  .I1(mux_o_2752),
  .S0(rad[6])
);
MUX2 mux_inst_2774 (
  .O(mux_o_2774),
  .I0(mux_o_2753),
  .I1(mux_o_2754),
  .S0(rad[6])
);
MUX2 mux_inst_2775 (
  .O(mux_o_2775),
  .I0(mux_o_2755),
  .I1(mux_o_2756),
  .S0(rad[6])
);
MUX2 mux_inst_2776 (
  .O(mux_o_2776),
  .I0(mux_o_2757),
  .I1(mux_o_2758),
  .S0(rad[6])
);
MUX2 mux_inst_2777 (
  .O(mux_o_2777),
  .I0(mux_o_2759),
  .I1(mux_o_2760),
  .S0(rad[6])
);
MUX2 mux_inst_2778 (
  .O(mux_o_2778),
  .I0(mux_o_2761),
  .I1(mux_o_2762),
  .S0(rad[6])
);
MUX2 mux_inst_2779 (
  .O(mux_o_2779),
  .I0(mux_o_2763),
  .I1(mux_o_2764),
  .S0(rad[7])
);
MUX2 mux_inst_2780 (
  .O(mux_o_2780),
  .I0(mux_o_2765),
  .I1(mux_o_2766),
  .S0(rad[7])
);
MUX2 mux_inst_2781 (
  .O(mux_o_2781),
  .I0(mux_o_2767),
  .I1(mux_o_2768),
  .S0(rad[7])
);
MUX2 mux_inst_2782 (
  .O(mux_o_2782),
  .I0(mux_o_2769),
  .I1(mux_o_2770),
  .S0(rad[7])
);
MUX2 mux_inst_2783 (
  .O(mux_o_2783),
  .I0(mux_o_2771),
  .I1(mux_o_2772),
  .S0(rad[7])
);
MUX2 mux_inst_2784 (
  .O(mux_o_2784),
  .I0(mux_o_2773),
  .I1(mux_o_2774),
  .S0(rad[7])
);
MUX2 mux_inst_2785 (
  .O(mux_o_2785),
  .I0(mux_o_2775),
  .I1(mux_o_2776),
  .S0(rad[7])
);
MUX2 mux_inst_2786 (
  .O(mux_o_2786),
  .I0(mux_o_2777),
  .I1(mux_o_2778),
  .S0(rad[7])
);
MUX2 mux_inst_2787 (
  .O(mux_o_2787),
  .I0(mux_o_2779),
  .I1(mux_o_2780),
  .S0(rad[8])
);
MUX2 mux_inst_2788 (
  .O(mux_o_2788),
  .I0(mux_o_2781),
  .I1(mux_o_2782),
  .S0(rad[8])
);
MUX2 mux_inst_2789 (
  .O(mux_o_2789),
  .I0(mux_o_2783),
  .I1(mux_o_2784),
  .S0(rad[8])
);
MUX2 mux_inst_2790 (
  .O(mux_o_2790),
  .I0(mux_o_2785),
  .I1(mux_o_2786),
  .S0(rad[8])
);
MUX2 mux_inst_2791 (
  .O(mux_o_2791),
  .I0(mux_o_2787),
  .I1(mux_o_2788),
  .S0(rad[9])
);
MUX2 mux_inst_2792 (
  .O(mux_o_2792),
  .I0(mux_o_2789),
  .I1(mux_o_2790),
  .S0(rad[9])
);
MUX2 mux_inst_2793 (
  .O(dout[21]),
  .I0(mux_o_2791),
  .I1(mux_o_2792),
  .S0(rad[10])
);
MUX2 mux_inst_2794 (
  .O(mux_o_2794),
  .I0(ram16sdp_inst_5_dout[22]),
  .I1(ram16sdp_inst_13_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2795 (
  .O(mux_o_2795),
  .I0(ram16sdp_inst_21_dout[22]),
  .I1(ram16sdp_inst_29_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2796 (
  .O(mux_o_2796),
  .I0(ram16sdp_inst_37_dout[22]),
  .I1(ram16sdp_inst_45_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2797 (
  .O(mux_o_2797),
  .I0(ram16sdp_inst_53_dout[22]),
  .I1(ram16sdp_inst_61_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2798 (
  .O(mux_o_2798),
  .I0(ram16sdp_inst_69_dout[22]),
  .I1(ram16sdp_inst_77_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2799 (
  .O(mux_o_2799),
  .I0(ram16sdp_inst_85_dout[22]),
  .I1(ram16sdp_inst_93_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2800 (
  .O(mux_o_2800),
  .I0(ram16sdp_inst_101_dout[22]),
  .I1(ram16sdp_inst_109_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2801 (
  .O(mux_o_2801),
  .I0(ram16sdp_inst_117_dout[22]),
  .I1(ram16sdp_inst_125_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2802 (
  .O(mux_o_2802),
  .I0(ram16sdp_inst_133_dout[22]),
  .I1(ram16sdp_inst_141_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2803 (
  .O(mux_o_2803),
  .I0(ram16sdp_inst_149_dout[22]),
  .I1(ram16sdp_inst_157_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2804 (
  .O(mux_o_2804),
  .I0(ram16sdp_inst_165_dout[22]),
  .I1(ram16sdp_inst_173_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2805 (
  .O(mux_o_2805),
  .I0(ram16sdp_inst_181_dout[22]),
  .I1(ram16sdp_inst_189_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2806 (
  .O(mux_o_2806),
  .I0(ram16sdp_inst_197_dout[22]),
  .I1(ram16sdp_inst_205_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2807 (
  .O(mux_o_2807),
  .I0(ram16sdp_inst_213_dout[22]),
  .I1(ram16sdp_inst_221_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2808 (
  .O(mux_o_2808),
  .I0(ram16sdp_inst_229_dout[22]),
  .I1(ram16sdp_inst_237_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2809 (
  .O(mux_o_2809),
  .I0(ram16sdp_inst_245_dout[22]),
  .I1(ram16sdp_inst_253_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2810 (
  .O(mux_o_2810),
  .I0(ram16sdp_inst_261_dout[22]),
  .I1(ram16sdp_inst_269_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2811 (
  .O(mux_o_2811),
  .I0(ram16sdp_inst_277_dout[22]),
  .I1(ram16sdp_inst_285_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2812 (
  .O(mux_o_2812),
  .I0(ram16sdp_inst_293_dout[22]),
  .I1(ram16sdp_inst_301_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2813 (
  .O(mux_o_2813),
  .I0(ram16sdp_inst_309_dout[22]),
  .I1(ram16sdp_inst_317_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2814 (
  .O(mux_o_2814),
  .I0(ram16sdp_inst_325_dout[22]),
  .I1(ram16sdp_inst_333_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2815 (
  .O(mux_o_2815),
  .I0(ram16sdp_inst_341_dout[22]),
  .I1(ram16sdp_inst_349_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2816 (
  .O(mux_o_2816),
  .I0(ram16sdp_inst_357_dout[22]),
  .I1(ram16sdp_inst_365_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2817 (
  .O(mux_o_2817),
  .I0(ram16sdp_inst_373_dout[22]),
  .I1(ram16sdp_inst_381_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2818 (
  .O(mux_o_2818),
  .I0(ram16sdp_inst_389_dout[22]),
  .I1(ram16sdp_inst_397_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2819 (
  .O(mux_o_2819),
  .I0(ram16sdp_inst_405_dout[22]),
  .I1(ram16sdp_inst_413_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2820 (
  .O(mux_o_2820),
  .I0(ram16sdp_inst_421_dout[22]),
  .I1(ram16sdp_inst_429_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2821 (
  .O(mux_o_2821),
  .I0(ram16sdp_inst_437_dout[22]),
  .I1(ram16sdp_inst_445_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2822 (
  .O(mux_o_2822),
  .I0(ram16sdp_inst_453_dout[22]),
  .I1(ram16sdp_inst_461_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2823 (
  .O(mux_o_2823),
  .I0(ram16sdp_inst_469_dout[22]),
  .I1(ram16sdp_inst_477_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2824 (
  .O(mux_o_2824),
  .I0(ram16sdp_inst_485_dout[22]),
  .I1(ram16sdp_inst_493_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2825 (
  .O(mux_o_2825),
  .I0(ram16sdp_inst_501_dout[22]),
  .I1(ram16sdp_inst_509_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2826 (
  .O(mux_o_2826),
  .I0(ram16sdp_inst_517_dout[22]),
  .I1(ram16sdp_inst_525_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2827 (
  .O(mux_o_2827),
  .I0(ram16sdp_inst_533_dout[22]),
  .I1(ram16sdp_inst_541_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2828 (
  .O(mux_o_2828),
  .I0(ram16sdp_inst_549_dout[22]),
  .I1(ram16sdp_inst_557_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2829 (
  .O(mux_o_2829),
  .I0(ram16sdp_inst_565_dout[22]),
  .I1(ram16sdp_inst_573_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2830 (
  .O(mux_o_2830),
  .I0(ram16sdp_inst_581_dout[22]),
  .I1(ram16sdp_inst_589_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2831 (
  .O(mux_o_2831),
  .I0(ram16sdp_inst_597_dout[22]),
  .I1(ram16sdp_inst_605_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2832 (
  .O(mux_o_2832),
  .I0(ram16sdp_inst_613_dout[22]),
  .I1(ram16sdp_inst_621_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2833 (
  .O(mux_o_2833),
  .I0(ram16sdp_inst_629_dout[22]),
  .I1(ram16sdp_inst_637_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2834 (
  .O(mux_o_2834),
  .I0(ram16sdp_inst_645_dout[22]),
  .I1(ram16sdp_inst_653_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2835 (
  .O(mux_o_2835),
  .I0(ram16sdp_inst_661_dout[22]),
  .I1(ram16sdp_inst_669_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2836 (
  .O(mux_o_2836),
  .I0(ram16sdp_inst_677_dout[22]),
  .I1(ram16sdp_inst_685_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2837 (
  .O(mux_o_2837),
  .I0(ram16sdp_inst_693_dout[22]),
  .I1(ram16sdp_inst_701_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2838 (
  .O(mux_o_2838),
  .I0(ram16sdp_inst_709_dout[22]),
  .I1(ram16sdp_inst_717_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2839 (
  .O(mux_o_2839),
  .I0(ram16sdp_inst_725_dout[22]),
  .I1(ram16sdp_inst_733_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2840 (
  .O(mux_o_2840),
  .I0(ram16sdp_inst_741_dout[22]),
  .I1(ram16sdp_inst_749_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2841 (
  .O(mux_o_2841),
  .I0(ram16sdp_inst_757_dout[22]),
  .I1(ram16sdp_inst_765_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2842 (
  .O(mux_o_2842),
  .I0(ram16sdp_inst_773_dout[22]),
  .I1(ram16sdp_inst_781_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2843 (
  .O(mux_o_2843),
  .I0(ram16sdp_inst_789_dout[22]),
  .I1(ram16sdp_inst_797_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2844 (
  .O(mux_o_2844),
  .I0(ram16sdp_inst_805_dout[22]),
  .I1(ram16sdp_inst_813_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2845 (
  .O(mux_o_2845),
  .I0(ram16sdp_inst_821_dout[22]),
  .I1(ram16sdp_inst_829_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2846 (
  .O(mux_o_2846),
  .I0(ram16sdp_inst_837_dout[22]),
  .I1(ram16sdp_inst_845_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2847 (
  .O(mux_o_2847),
  .I0(ram16sdp_inst_853_dout[22]),
  .I1(ram16sdp_inst_861_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2848 (
  .O(mux_o_2848),
  .I0(ram16sdp_inst_869_dout[22]),
  .I1(ram16sdp_inst_877_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2849 (
  .O(mux_o_2849),
  .I0(ram16sdp_inst_885_dout[22]),
  .I1(ram16sdp_inst_893_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2850 (
  .O(mux_o_2850),
  .I0(ram16sdp_inst_901_dout[22]),
  .I1(ram16sdp_inst_909_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2851 (
  .O(mux_o_2851),
  .I0(ram16sdp_inst_917_dout[22]),
  .I1(ram16sdp_inst_925_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2852 (
  .O(mux_o_2852),
  .I0(ram16sdp_inst_933_dout[22]),
  .I1(ram16sdp_inst_941_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2853 (
  .O(mux_o_2853),
  .I0(ram16sdp_inst_949_dout[22]),
  .I1(ram16sdp_inst_957_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2854 (
  .O(mux_o_2854),
  .I0(ram16sdp_inst_965_dout[22]),
  .I1(ram16sdp_inst_973_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2855 (
  .O(mux_o_2855),
  .I0(ram16sdp_inst_981_dout[22]),
  .I1(ram16sdp_inst_989_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2856 (
  .O(mux_o_2856),
  .I0(ram16sdp_inst_997_dout[22]),
  .I1(ram16sdp_inst_1005_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2857 (
  .O(mux_o_2857),
  .I0(ram16sdp_inst_1013_dout[22]),
  .I1(ram16sdp_inst_1021_dout[22]),
  .S0(rad[4])
);
MUX2 mux_inst_2858 (
  .O(mux_o_2858),
  .I0(mux_o_2794),
  .I1(mux_o_2795),
  .S0(rad[5])
);
MUX2 mux_inst_2859 (
  .O(mux_o_2859),
  .I0(mux_o_2796),
  .I1(mux_o_2797),
  .S0(rad[5])
);
MUX2 mux_inst_2860 (
  .O(mux_o_2860),
  .I0(mux_o_2798),
  .I1(mux_o_2799),
  .S0(rad[5])
);
MUX2 mux_inst_2861 (
  .O(mux_o_2861),
  .I0(mux_o_2800),
  .I1(mux_o_2801),
  .S0(rad[5])
);
MUX2 mux_inst_2862 (
  .O(mux_o_2862),
  .I0(mux_o_2802),
  .I1(mux_o_2803),
  .S0(rad[5])
);
MUX2 mux_inst_2863 (
  .O(mux_o_2863),
  .I0(mux_o_2804),
  .I1(mux_o_2805),
  .S0(rad[5])
);
MUX2 mux_inst_2864 (
  .O(mux_o_2864),
  .I0(mux_o_2806),
  .I1(mux_o_2807),
  .S0(rad[5])
);
MUX2 mux_inst_2865 (
  .O(mux_o_2865),
  .I0(mux_o_2808),
  .I1(mux_o_2809),
  .S0(rad[5])
);
MUX2 mux_inst_2866 (
  .O(mux_o_2866),
  .I0(mux_o_2810),
  .I1(mux_o_2811),
  .S0(rad[5])
);
MUX2 mux_inst_2867 (
  .O(mux_o_2867),
  .I0(mux_o_2812),
  .I1(mux_o_2813),
  .S0(rad[5])
);
MUX2 mux_inst_2868 (
  .O(mux_o_2868),
  .I0(mux_o_2814),
  .I1(mux_o_2815),
  .S0(rad[5])
);
MUX2 mux_inst_2869 (
  .O(mux_o_2869),
  .I0(mux_o_2816),
  .I1(mux_o_2817),
  .S0(rad[5])
);
MUX2 mux_inst_2870 (
  .O(mux_o_2870),
  .I0(mux_o_2818),
  .I1(mux_o_2819),
  .S0(rad[5])
);
MUX2 mux_inst_2871 (
  .O(mux_o_2871),
  .I0(mux_o_2820),
  .I1(mux_o_2821),
  .S0(rad[5])
);
MUX2 mux_inst_2872 (
  .O(mux_o_2872),
  .I0(mux_o_2822),
  .I1(mux_o_2823),
  .S0(rad[5])
);
MUX2 mux_inst_2873 (
  .O(mux_o_2873),
  .I0(mux_o_2824),
  .I1(mux_o_2825),
  .S0(rad[5])
);
MUX2 mux_inst_2874 (
  .O(mux_o_2874),
  .I0(mux_o_2826),
  .I1(mux_o_2827),
  .S0(rad[5])
);
MUX2 mux_inst_2875 (
  .O(mux_o_2875),
  .I0(mux_o_2828),
  .I1(mux_o_2829),
  .S0(rad[5])
);
MUX2 mux_inst_2876 (
  .O(mux_o_2876),
  .I0(mux_o_2830),
  .I1(mux_o_2831),
  .S0(rad[5])
);
MUX2 mux_inst_2877 (
  .O(mux_o_2877),
  .I0(mux_o_2832),
  .I1(mux_o_2833),
  .S0(rad[5])
);
MUX2 mux_inst_2878 (
  .O(mux_o_2878),
  .I0(mux_o_2834),
  .I1(mux_o_2835),
  .S0(rad[5])
);
MUX2 mux_inst_2879 (
  .O(mux_o_2879),
  .I0(mux_o_2836),
  .I1(mux_o_2837),
  .S0(rad[5])
);
MUX2 mux_inst_2880 (
  .O(mux_o_2880),
  .I0(mux_o_2838),
  .I1(mux_o_2839),
  .S0(rad[5])
);
MUX2 mux_inst_2881 (
  .O(mux_o_2881),
  .I0(mux_o_2840),
  .I1(mux_o_2841),
  .S0(rad[5])
);
MUX2 mux_inst_2882 (
  .O(mux_o_2882),
  .I0(mux_o_2842),
  .I1(mux_o_2843),
  .S0(rad[5])
);
MUX2 mux_inst_2883 (
  .O(mux_o_2883),
  .I0(mux_o_2844),
  .I1(mux_o_2845),
  .S0(rad[5])
);
MUX2 mux_inst_2884 (
  .O(mux_o_2884),
  .I0(mux_o_2846),
  .I1(mux_o_2847),
  .S0(rad[5])
);
MUX2 mux_inst_2885 (
  .O(mux_o_2885),
  .I0(mux_o_2848),
  .I1(mux_o_2849),
  .S0(rad[5])
);
MUX2 mux_inst_2886 (
  .O(mux_o_2886),
  .I0(mux_o_2850),
  .I1(mux_o_2851),
  .S0(rad[5])
);
MUX2 mux_inst_2887 (
  .O(mux_o_2887),
  .I0(mux_o_2852),
  .I1(mux_o_2853),
  .S0(rad[5])
);
MUX2 mux_inst_2888 (
  .O(mux_o_2888),
  .I0(mux_o_2854),
  .I1(mux_o_2855),
  .S0(rad[5])
);
MUX2 mux_inst_2889 (
  .O(mux_o_2889),
  .I0(mux_o_2856),
  .I1(mux_o_2857),
  .S0(rad[5])
);
MUX2 mux_inst_2890 (
  .O(mux_o_2890),
  .I0(mux_o_2858),
  .I1(mux_o_2859),
  .S0(rad[6])
);
MUX2 mux_inst_2891 (
  .O(mux_o_2891),
  .I0(mux_o_2860),
  .I1(mux_o_2861),
  .S0(rad[6])
);
MUX2 mux_inst_2892 (
  .O(mux_o_2892),
  .I0(mux_o_2862),
  .I1(mux_o_2863),
  .S0(rad[6])
);
MUX2 mux_inst_2893 (
  .O(mux_o_2893),
  .I0(mux_o_2864),
  .I1(mux_o_2865),
  .S0(rad[6])
);
MUX2 mux_inst_2894 (
  .O(mux_o_2894),
  .I0(mux_o_2866),
  .I1(mux_o_2867),
  .S0(rad[6])
);
MUX2 mux_inst_2895 (
  .O(mux_o_2895),
  .I0(mux_o_2868),
  .I1(mux_o_2869),
  .S0(rad[6])
);
MUX2 mux_inst_2896 (
  .O(mux_o_2896),
  .I0(mux_o_2870),
  .I1(mux_o_2871),
  .S0(rad[6])
);
MUX2 mux_inst_2897 (
  .O(mux_o_2897),
  .I0(mux_o_2872),
  .I1(mux_o_2873),
  .S0(rad[6])
);
MUX2 mux_inst_2898 (
  .O(mux_o_2898),
  .I0(mux_o_2874),
  .I1(mux_o_2875),
  .S0(rad[6])
);
MUX2 mux_inst_2899 (
  .O(mux_o_2899),
  .I0(mux_o_2876),
  .I1(mux_o_2877),
  .S0(rad[6])
);
MUX2 mux_inst_2900 (
  .O(mux_o_2900),
  .I0(mux_o_2878),
  .I1(mux_o_2879),
  .S0(rad[6])
);
MUX2 mux_inst_2901 (
  .O(mux_o_2901),
  .I0(mux_o_2880),
  .I1(mux_o_2881),
  .S0(rad[6])
);
MUX2 mux_inst_2902 (
  .O(mux_o_2902),
  .I0(mux_o_2882),
  .I1(mux_o_2883),
  .S0(rad[6])
);
MUX2 mux_inst_2903 (
  .O(mux_o_2903),
  .I0(mux_o_2884),
  .I1(mux_o_2885),
  .S0(rad[6])
);
MUX2 mux_inst_2904 (
  .O(mux_o_2904),
  .I0(mux_o_2886),
  .I1(mux_o_2887),
  .S0(rad[6])
);
MUX2 mux_inst_2905 (
  .O(mux_o_2905),
  .I0(mux_o_2888),
  .I1(mux_o_2889),
  .S0(rad[6])
);
MUX2 mux_inst_2906 (
  .O(mux_o_2906),
  .I0(mux_o_2890),
  .I1(mux_o_2891),
  .S0(rad[7])
);
MUX2 mux_inst_2907 (
  .O(mux_o_2907),
  .I0(mux_o_2892),
  .I1(mux_o_2893),
  .S0(rad[7])
);
MUX2 mux_inst_2908 (
  .O(mux_o_2908),
  .I0(mux_o_2894),
  .I1(mux_o_2895),
  .S0(rad[7])
);
MUX2 mux_inst_2909 (
  .O(mux_o_2909),
  .I0(mux_o_2896),
  .I1(mux_o_2897),
  .S0(rad[7])
);
MUX2 mux_inst_2910 (
  .O(mux_o_2910),
  .I0(mux_o_2898),
  .I1(mux_o_2899),
  .S0(rad[7])
);
MUX2 mux_inst_2911 (
  .O(mux_o_2911),
  .I0(mux_o_2900),
  .I1(mux_o_2901),
  .S0(rad[7])
);
MUX2 mux_inst_2912 (
  .O(mux_o_2912),
  .I0(mux_o_2902),
  .I1(mux_o_2903),
  .S0(rad[7])
);
MUX2 mux_inst_2913 (
  .O(mux_o_2913),
  .I0(mux_o_2904),
  .I1(mux_o_2905),
  .S0(rad[7])
);
MUX2 mux_inst_2914 (
  .O(mux_o_2914),
  .I0(mux_o_2906),
  .I1(mux_o_2907),
  .S0(rad[8])
);
MUX2 mux_inst_2915 (
  .O(mux_o_2915),
  .I0(mux_o_2908),
  .I1(mux_o_2909),
  .S0(rad[8])
);
MUX2 mux_inst_2916 (
  .O(mux_o_2916),
  .I0(mux_o_2910),
  .I1(mux_o_2911),
  .S0(rad[8])
);
MUX2 mux_inst_2917 (
  .O(mux_o_2917),
  .I0(mux_o_2912),
  .I1(mux_o_2913),
  .S0(rad[8])
);
MUX2 mux_inst_2918 (
  .O(mux_o_2918),
  .I0(mux_o_2914),
  .I1(mux_o_2915),
  .S0(rad[9])
);
MUX2 mux_inst_2919 (
  .O(mux_o_2919),
  .I0(mux_o_2916),
  .I1(mux_o_2917),
  .S0(rad[9])
);
MUX2 mux_inst_2920 (
  .O(dout[22]),
  .I0(mux_o_2918),
  .I1(mux_o_2919),
  .S0(rad[10])
);
MUX2 mux_inst_2921 (
  .O(mux_o_2921),
  .I0(ram16sdp_inst_5_dout[23]),
  .I1(ram16sdp_inst_13_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2922 (
  .O(mux_o_2922),
  .I0(ram16sdp_inst_21_dout[23]),
  .I1(ram16sdp_inst_29_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2923 (
  .O(mux_o_2923),
  .I0(ram16sdp_inst_37_dout[23]),
  .I1(ram16sdp_inst_45_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2924 (
  .O(mux_o_2924),
  .I0(ram16sdp_inst_53_dout[23]),
  .I1(ram16sdp_inst_61_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2925 (
  .O(mux_o_2925),
  .I0(ram16sdp_inst_69_dout[23]),
  .I1(ram16sdp_inst_77_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2926 (
  .O(mux_o_2926),
  .I0(ram16sdp_inst_85_dout[23]),
  .I1(ram16sdp_inst_93_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2927 (
  .O(mux_o_2927),
  .I0(ram16sdp_inst_101_dout[23]),
  .I1(ram16sdp_inst_109_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2928 (
  .O(mux_o_2928),
  .I0(ram16sdp_inst_117_dout[23]),
  .I1(ram16sdp_inst_125_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2929 (
  .O(mux_o_2929),
  .I0(ram16sdp_inst_133_dout[23]),
  .I1(ram16sdp_inst_141_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2930 (
  .O(mux_o_2930),
  .I0(ram16sdp_inst_149_dout[23]),
  .I1(ram16sdp_inst_157_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2931 (
  .O(mux_o_2931),
  .I0(ram16sdp_inst_165_dout[23]),
  .I1(ram16sdp_inst_173_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2932 (
  .O(mux_o_2932),
  .I0(ram16sdp_inst_181_dout[23]),
  .I1(ram16sdp_inst_189_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2933 (
  .O(mux_o_2933),
  .I0(ram16sdp_inst_197_dout[23]),
  .I1(ram16sdp_inst_205_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2934 (
  .O(mux_o_2934),
  .I0(ram16sdp_inst_213_dout[23]),
  .I1(ram16sdp_inst_221_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2935 (
  .O(mux_o_2935),
  .I0(ram16sdp_inst_229_dout[23]),
  .I1(ram16sdp_inst_237_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2936 (
  .O(mux_o_2936),
  .I0(ram16sdp_inst_245_dout[23]),
  .I1(ram16sdp_inst_253_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2937 (
  .O(mux_o_2937),
  .I0(ram16sdp_inst_261_dout[23]),
  .I1(ram16sdp_inst_269_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2938 (
  .O(mux_o_2938),
  .I0(ram16sdp_inst_277_dout[23]),
  .I1(ram16sdp_inst_285_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2939 (
  .O(mux_o_2939),
  .I0(ram16sdp_inst_293_dout[23]),
  .I1(ram16sdp_inst_301_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2940 (
  .O(mux_o_2940),
  .I0(ram16sdp_inst_309_dout[23]),
  .I1(ram16sdp_inst_317_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2941 (
  .O(mux_o_2941),
  .I0(ram16sdp_inst_325_dout[23]),
  .I1(ram16sdp_inst_333_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2942 (
  .O(mux_o_2942),
  .I0(ram16sdp_inst_341_dout[23]),
  .I1(ram16sdp_inst_349_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2943 (
  .O(mux_o_2943),
  .I0(ram16sdp_inst_357_dout[23]),
  .I1(ram16sdp_inst_365_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2944 (
  .O(mux_o_2944),
  .I0(ram16sdp_inst_373_dout[23]),
  .I1(ram16sdp_inst_381_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2945 (
  .O(mux_o_2945),
  .I0(ram16sdp_inst_389_dout[23]),
  .I1(ram16sdp_inst_397_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2946 (
  .O(mux_o_2946),
  .I0(ram16sdp_inst_405_dout[23]),
  .I1(ram16sdp_inst_413_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2947 (
  .O(mux_o_2947),
  .I0(ram16sdp_inst_421_dout[23]),
  .I1(ram16sdp_inst_429_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2948 (
  .O(mux_o_2948),
  .I0(ram16sdp_inst_437_dout[23]),
  .I1(ram16sdp_inst_445_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2949 (
  .O(mux_o_2949),
  .I0(ram16sdp_inst_453_dout[23]),
  .I1(ram16sdp_inst_461_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2950 (
  .O(mux_o_2950),
  .I0(ram16sdp_inst_469_dout[23]),
  .I1(ram16sdp_inst_477_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2951 (
  .O(mux_o_2951),
  .I0(ram16sdp_inst_485_dout[23]),
  .I1(ram16sdp_inst_493_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2952 (
  .O(mux_o_2952),
  .I0(ram16sdp_inst_501_dout[23]),
  .I1(ram16sdp_inst_509_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2953 (
  .O(mux_o_2953),
  .I0(ram16sdp_inst_517_dout[23]),
  .I1(ram16sdp_inst_525_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2954 (
  .O(mux_o_2954),
  .I0(ram16sdp_inst_533_dout[23]),
  .I1(ram16sdp_inst_541_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2955 (
  .O(mux_o_2955),
  .I0(ram16sdp_inst_549_dout[23]),
  .I1(ram16sdp_inst_557_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2956 (
  .O(mux_o_2956),
  .I0(ram16sdp_inst_565_dout[23]),
  .I1(ram16sdp_inst_573_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2957 (
  .O(mux_o_2957),
  .I0(ram16sdp_inst_581_dout[23]),
  .I1(ram16sdp_inst_589_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2958 (
  .O(mux_o_2958),
  .I0(ram16sdp_inst_597_dout[23]),
  .I1(ram16sdp_inst_605_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2959 (
  .O(mux_o_2959),
  .I0(ram16sdp_inst_613_dout[23]),
  .I1(ram16sdp_inst_621_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2960 (
  .O(mux_o_2960),
  .I0(ram16sdp_inst_629_dout[23]),
  .I1(ram16sdp_inst_637_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2961 (
  .O(mux_o_2961),
  .I0(ram16sdp_inst_645_dout[23]),
  .I1(ram16sdp_inst_653_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2962 (
  .O(mux_o_2962),
  .I0(ram16sdp_inst_661_dout[23]),
  .I1(ram16sdp_inst_669_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2963 (
  .O(mux_o_2963),
  .I0(ram16sdp_inst_677_dout[23]),
  .I1(ram16sdp_inst_685_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2964 (
  .O(mux_o_2964),
  .I0(ram16sdp_inst_693_dout[23]),
  .I1(ram16sdp_inst_701_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2965 (
  .O(mux_o_2965),
  .I0(ram16sdp_inst_709_dout[23]),
  .I1(ram16sdp_inst_717_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2966 (
  .O(mux_o_2966),
  .I0(ram16sdp_inst_725_dout[23]),
  .I1(ram16sdp_inst_733_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2967 (
  .O(mux_o_2967),
  .I0(ram16sdp_inst_741_dout[23]),
  .I1(ram16sdp_inst_749_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2968 (
  .O(mux_o_2968),
  .I0(ram16sdp_inst_757_dout[23]),
  .I1(ram16sdp_inst_765_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2969 (
  .O(mux_o_2969),
  .I0(ram16sdp_inst_773_dout[23]),
  .I1(ram16sdp_inst_781_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2970 (
  .O(mux_o_2970),
  .I0(ram16sdp_inst_789_dout[23]),
  .I1(ram16sdp_inst_797_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2971 (
  .O(mux_o_2971),
  .I0(ram16sdp_inst_805_dout[23]),
  .I1(ram16sdp_inst_813_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2972 (
  .O(mux_o_2972),
  .I0(ram16sdp_inst_821_dout[23]),
  .I1(ram16sdp_inst_829_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2973 (
  .O(mux_o_2973),
  .I0(ram16sdp_inst_837_dout[23]),
  .I1(ram16sdp_inst_845_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2974 (
  .O(mux_o_2974),
  .I0(ram16sdp_inst_853_dout[23]),
  .I1(ram16sdp_inst_861_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2975 (
  .O(mux_o_2975),
  .I0(ram16sdp_inst_869_dout[23]),
  .I1(ram16sdp_inst_877_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2976 (
  .O(mux_o_2976),
  .I0(ram16sdp_inst_885_dout[23]),
  .I1(ram16sdp_inst_893_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2977 (
  .O(mux_o_2977),
  .I0(ram16sdp_inst_901_dout[23]),
  .I1(ram16sdp_inst_909_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2978 (
  .O(mux_o_2978),
  .I0(ram16sdp_inst_917_dout[23]),
  .I1(ram16sdp_inst_925_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2979 (
  .O(mux_o_2979),
  .I0(ram16sdp_inst_933_dout[23]),
  .I1(ram16sdp_inst_941_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2980 (
  .O(mux_o_2980),
  .I0(ram16sdp_inst_949_dout[23]),
  .I1(ram16sdp_inst_957_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2981 (
  .O(mux_o_2981),
  .I0(ram16sdp_inst_965_dout[23]),
  .I1(ram16sdp_inst_973_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2982 (
  .O(mux_o_2982),
  .I0(ram16sdp_inst_981_dout[23]),
  .I1(ram16sdp_inst_989_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2983 (
  .O(mux_o_2983),
  .I0(ram16sdp_inst_997_dout[23]),
  .I1(ram16sdp_inst_1005_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2984 (
  .O(mux_o_2984),
  .I0(ram16sdp_inst_1013_dout[23]),
  .I1(ram16sdp_inst_1021_dout[23]),
  .S0(rad[4])
);
MUX2 mux_inst_2985 (
  .O(mux_o_2985),
  .I0(mux_o_2921),
  .I1(mux_o_2922),
  .S0(rad[5])
);
MUX2 mux_inst_2986 (
  .O(mux_o_2986),
  .I0(mux_o_2923),
  .I1(mux_o_2924),
  .S0(rad[5])
);
MUX2 mux_inst_2987 (
  .O(mux_o_2987),
  .I0(mux_o_2925),
  .I1(mux_o_2926),
  .S0(rad[5])
);
MUX2 mux_inst_2988 (
  .O(mux_o_2988),
  .I0(mux_o_2927),
  .I1(mux_o_2928),
  .S0(rad[5])
);
MUX2 mux_inst_2989 (
  .O(mux_o_2989),
  .I0(mux_o_2929),
  .I1(mux_o_2930),
  .S0(rad[5])
);
MUX2 mux_inst_2990 (
  .O(mux_o_2990),
  .I0(mux_o_2931),
  .I1(mux_o_2932),
  .S0(rad[5])
);
MUX2 mux_inst_2991 (
  .O(mux_o_2991),
  .I0(mux_o_2933),
  .I1(mux_o_2934),
  .S0(rad[5])
);
MUX2 mux_inst_2992 (
  .O(mux_o_2992),
  .I0(mux_o_2935),
  .I1(mux_o_2936),
  .S0(rad[5])
);
MUX2 mux_inst_2993 (
  .O(mux_o_2993),
  .I0(mux_o_2937),
  .I1(mux_o_2938),
  .S0(rad[5])
);
MUX2 mux_inst_2994 (
  .O(mux_o_2994),
  .I0(mux_o_2939),
  .I1(mux_o_2940),
  .S0(rad[5])
);
MUX2 mux_inst_2995 (
  .O(mux_o_2995),
  .I0(mux_o_2941),
  .I1(mux_o_2942),
  .S0(rad[5])
);
MUX2 mux_inst_2996 (
  .O(mux_o_2996),
  .I0(mux_o_2943),
  .I1(mux_o_2944),
  .S0(rad[5])
);
MUX2 mux_inst_2997 (
  .O(mux_o_2997),
  .I0(mux_o_2945),
  .I1(mux_o_2946),
  .S0(rad[5])
);
MUX2 mux_inst_2998 (
  .O(mux_o_2998),
  .I0(mux_o_2947),
  .I1(mux_o_2948),
  .S0(rad[5])
);
MUX2 mux_inst_2999 (
  .O(mux_o_2999),
  .I0(mux_o_2949),
  .I1(mux_o_2950),
  .S0(rad[5])
);
MUX2 mux_inst_3000 (
  .O(mux_o_3000),
  .I0(mux_o_2951),
  .I1(mux_o_2952),
  .S0(rad[5])
);
MUX2 mux_inst_3001 (
  .O(mux_o_3001),
  .I0(mux_o_2953),
  .I1(mux_o_2954),
  .S0(rad[5])
);
MUX2 mux_inst_3002 (
  .O(mux_o_3002),
  .I0(mux_o_2955),
  .I1(mux_o_2956),
  .S0(rad[5])
);
MUX2 mux_inst_3003 (
  .O(mux_o_3003),
  .I0(mux_o_2957),
  .I1(mux_o_2958),
  .S0(rad[5])
);
MUX2 mux_inst_3004 (
  .O(mux_o_3004),
  .I0(mux_o_2959),
  .I1(mux_o_2960),
  .S0(rad[5])
);
MUX2 mux_inst_3005 (
  .O(mux_o_3005),
  .I0(mux_o_2961),
  .I1(mux_o_2962),
  .S0(rad[5])
);
MUX2 mux_inst_3006 (
  .O(mux_o_3006),
  .I0(mux_o_2963),
  .I1(mux_o_2964),
  .S0(rad[5])
);
MUX2 mux_inst_3007 (
  .O(mux_o_3007),
  .I0(mux_o_2965),
  .I1(mux_o_2966),
  .S0(rad[5])
);
MUX2 mux_inst_3008 (
  .O(mux_o_3008),
  .I0(mux_o_2967),
  .I1(mux_o_2968),
  .S0(rad[5])
);
MUX2 mux_inst_3009 (
  .O(mux_o_3009),
  .I0(mux_o_2969),
  .I1(mux_o_2970),
  .S0(rad[5])
);
MUX2 mux_inst_3010 (
  .O(mux_o_3010),
  .I0(mux_o_2971),
  .I1(mux_o_2972),
  .S0(rad[5])
);
MUX2 mux_inst_3011 (
  .O(mux_o_3011),
  .I0(mux_o_2973),
  .I1(mux_o_2974),
  .S0(rad[5])
);
MUX2 mux_inst_3012 (
  .O(mux_o_3012),
  .I0(mux_o_2975),
  .I1(mux_o_2976),
  .S0(rad[5])
);
MUX2 mux_inst_3013 (
  .O(mux_o_3013),
  .I0(mux_o_2977),
  .I1(mux_o_2978),
  .S0(rad[5])
);
MUX2 mux_inst_3014 (
  .O(mux_o_3014),
  .I0(mux_o_2979),
  .I1(mux_o_2980),
  .S0(rad[5])
);
MUX2 mux_inst_3015 (
  .O(mux_o_3015),
  .I0(mux_o_2981),
  .I1(mux_o_2982),
  .S0(rad[5])
);
MUX2 mux_inst_3016 (
  .O(mux_o_3016),
  .I0(mux_o_2983),
  .I1(mux_o_2984),
  .S0(rad[5])
);
MUX2 mux_inst_3017 (
  .O(mux_o_3017),
  .I0(mux_o_2985),
  .I1(mux_o_2986),
  .S0(rad[6])
);
MUX2 mux_inst_3018 (
  .O(mux_o_3018),
  .I0(mux_o_2987),
  .I1(mux_o_2988),
  .S0(rad[6])
);
MUX2 mux_inst_3019 (
  .O(mux_o_3019),
  .I0(mux_o_2989),
  .I1(mux_o_2990),
  .S0(rad[6])
);
MUX2 mux_inst_3020 (
  .O(mux_o_3020),
  .I0(mux_o_2991),
  .I1(mux_o_2992),
  .S0(rad[6])
);
MUX2 mux_inst_3021 (
  .O(mux_o_3021),
  .I0(mux_o_2993),
  .I1(mux_o_2994),
  .S0(rad[6])
);
MUX2 mux_inst_3022 (
  .O(mux_o_3022),
  .I0(mux_o_2995),
  .I1(mux_o_2996),
  .S0(rad[6])
);
MUX2 mux_inst_3023 (
  .O(mux_o_3023),
  .I0(mux_o_2997),
  .I1(mux_o_2998),
  .S0(rad[6])
);
MUX2 mux_inst_3024 (
  .O(mux_o_3024),
  .I0(mux_o_2999),
  .I1(mux_o_3000),
  .S0(rad[6])
);
MUX2 mux_inst_3025 (
  .O(mux_o_3025),
  .I0(mux_o_3001),
  .I1(mux_o_3002),
  .S0(rad[6])
);
MUX2 mux_inst_3026 (
  .O(mux_o_3026),
  .I0(mux_o_3003),
  .I1(mux_o_3004),
  .S0(rad[6])
);
MUX2 mux_inst_3027 (
  .O(mux_o_3027),
  .I0(mux_o_3005),
  .I1(mux_o_3006),
  .S0(rad[6])
);
MUX2 mux_inst_3028 (
  .O(mux_o_3028),
  .I0(mux_o_3007),
  .I1(mux_o_3008),
  .S0(rad[6])
);
MUX2 mux_inst_3029 (
  .O(mux_o_3029),
  .I0(mux_o_3009),
  .I1(mux_o_3010),
  .S0(rad[6])
);
MUX2 mux_inst_3030 (
  .O(mux_o_3030),
  .I0(mux_o_3011),
  .I1(mux_o_3012),
  .S0(rad[6])
);
MUX2 mux_inst_3031 (
  .O(mux_o_3031),
  .I0(mux_o_3013),
  .I1(mux_o_3014),
  .S0(rad[6])
);
MUX2 mux_inst_3032 (
  .O(mux_o_3032),
  .I0(mux_o_3015),
  .I1(mux_o_3016),
  .S0(rad[6])
);
MUX2 mux_inst_3033 (
  .O(mux_o_3033),
  .I0(mux_o_3017),
  .I1(mux_o_3018),
  .S0(rad[7])
);
MUX2 mux_inst_3034 (
  .O(mux_o_3034),
  .I0(mux_o_3019),
  .I1(mux_o_3020),
  .S0(rad[7])
);
MUX2 mux_inst_3035 (
  .O(mux_o_3035),
  .I0(mux_o_3021),
  .I1(mux_o_3022),
  .S0(rad[7])
);
MUX2 mux_inst_3036 (
  .O(mux_o_3036),
  .I0(mux_o_3023),
  .I1(mux_o_3024),
  .S0(rad[7])
);
MUX2 mux_inst_3037 (
  .O(mux_o_3037),
  .I0(mux_o_3025),
  .I1(mux_o_3026),
  .S0(rad[7])
);
MUX2 mux_inst_3038 (
  .O(mux_o_3038),
  .I0(mux_o_3027),
  .I1(mux_o_3028),
  .S0(rad[7])
);
MUX2 mux_inst_3039 (
  .O(mux_o_3039),
  .I0(mux_o_3029),
  .I1(mux_o_3030),
  .S0(rad[7])
);
MUX2 mux_inst_3040 (
  .O(mux_o_3040),
  .I0(mux_o_3031),
  .I1(mux_o_3032),
  .S0(rad[7])
);
MUX2 mux_inst_3041 (
  .O(mux_o_3041),
  .I0(mux_o_3033),
  .I1(mux_o_3034),
  .S0(rad[8])
);
MUX2 mux_inst_3042 (
  .O(mux_o_3042),
  .I0(mux_o_3035),
  .I1(mux_o_3036),
  .S0(rad[8])
);
MUX2 mux_inst_3043 (
  .O(mux_o_3043),
  .I0(mux_o_3037),
  .I1(mux_o_3038),
  .S0(rad[8])
);
MUX2 mux_inst_3044 (
  .O(mux_o_3044),
  .I0(mux_o_3039),
  .I1(mux_o_3040),
  .S0(rad[8])
);
MUX2 mux_inst_3045 (
  .O(mux_o_3045),
  .I0(mux_o_3041),
  .I1(mux_o_3042),
  .S0(rad[9])
);
MUX2 mux_inst_3046 (
  .O(mux_o_3046),
  .I0(mux_o_3043),
  .I1(mux_o_3044),
  .S0(rad[9])
);
MUX2 mux_inst_3047 (
  .O(dout[23]),
  .I0(mux_o_3045),
  .I1(mux_o_3046),
  .S0(rad[10])
);
MUX2 mux_inst_3048 (
  .O(mux_o_3048),
  .I0(ram16sdp_inst_6_dout[24]),
  .I1(ram16sdp_inst_14_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3049 (
  .O(mux_o_3049),
  .I0(ram16sdp_inst_22_dout[24]),
  .I1(ram16sdp_inst_30_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3050 (
  .O(mux_o_3050),
  .I0(ram16sdp_inst_38_dout[24]),
  .I1(ram16sdp_inst_46_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3051 (
  .O(mux_o_3051),
  .I0(ram16sdp_inst_54_dout[24]),
  .I1(ram16sdp_inst_62_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3052 (
  .O(mux_o_3052),
  .I0(ram16sdp_inst_70_dout[24]),
  .I1(ram16sdp_inst_78_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3053 (
  .O(mux_o_3053),
  .I0(ram16sdp_inst_86_dout[24]),
  .I1(ram16sdp_inst_94_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3054 (
  .O(mux_o_3054),
  .I0(ram16sdp_inst_102_dout[24]),
  .I1(ram16sdp_inst_110_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3055 (
  .O(mux_o_3055),
  .I0(ram16sdp_inst_118_dout[24]),
  .I1(ram16sdp_inst_126_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3056 (
  .O(mux_o_3056),
  .I0(ram16sdp_inst_134_dout[24]),
  .I1(ram16sdp_inst_142_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3057 (
  .O(mux_o_3057),
  .I0(ram16sdp_inst_150_dout[24]),
  .I1(ram16sdp_inst_158_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3058 (
  .O(mux_o_3058),
  .I0(ram16sdp_inst_166_dout[24]),
  .I1(ram16sdp_inst_174_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3059 (
  .O(mux_o_3059),
  .I0(ram16sdp_inst_182_dout[24]),
  .I1(ram16sdp_inst_190_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3060 (
  .O(mux_o_3060),
  .I0(ram16sdp_inst_198_dout[24]),
  .I1(ram16sdp_inst_206_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3061 (
  .O(mux_o_3061),
  .I0(ram16sdp_inst_214_dout[24]),
  .I1(ram16sdp_inst_222_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3062 (
  .O(mux_o_3062),
  .I0(ram16sdp_inst_230_dout[24]),
  .I1(ram16sdp_inst_238_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3063 (
  .O(mux_o_3063),
  .I0(ram16sdp_inst_246_dout[24]),
  .I1(ram16sdp_inst_254_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3064 (
  .O(mux_o_3064),
  .I0(ram16sdp_inst_262_dout[24]),
  .I1(ram16sdp_inst_270_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3065 (
  .O(mux_o_3065),
  .I0(ram16sdp_inst_278_dout[24]),
  .I1(ram16sdp_inst_286_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3066 (
  .O(mux_o_3066),
  .I0(ram16sdp_inst_294_dout[24]),
  .I1(ram16sdp_inst_302_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3067 (
  .O(mux_o_3067),
  .I0(ram16sdp_inst_310_dout[24]),
  .I1(ram16sdp_inst_318_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3068 (
  .O(mux_o_3068),
  .I0(ram16sdp_inst_326_dout[24]),
  .I1(ram16sdp_inst_334_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3069 (
  .O(mux_o_3069),
  .I0(ram16sdp_inst_342_dout[24]),
  .I1(ram16sdp_inst_350_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3070 (
  .O(mux_o_3070),
  .I0(ram16sdp_inst_358_dout[24]),
  .I1(ram16sdp_inst_366_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3071 (
  .O(mux_o_3071),
  .I0(ram16sdp_inst_374_dout[24]),
  .I1(ram16sdp_inst_382_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3072 (
  .O(mux_o_3072),
  .I0(ram16sdp_inst_390_dout[24]),
  .I1(ram16sdp_inst_398_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3073 (
  .O(mux_o_3073),
  .I0(ram16sdp_inst_406_dout[24]),
  .I1(ram16sdp_inst_414_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3074 (
  .O(mux_o_3074),
  .I0(ram16sdp_inst_422_dout[24]),
  .I1(ram16sdp_inst_430_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3075 (
  .O(mux_o_3075),
  .I0(ram16sdp_inst_438_dout[24]),
  .I1(ram16sdp_inst_446_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3076 (
  .O(mux_o_3076),
  .I0(ram16sdp_inst_454_dout[24]),
  .I1(ram16sdp_inst_462_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3077 (
  .O(mux_o_3077),
  .I0(ram16sdp_inst_470_dout[24]),
  .I1(ram16sdp_inst_478_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3078 (
  .O(mux_o_3078),
  .I0(ram16sdp_inst_486_dout[24]),
  .I1(ram16sdp_inst_494_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3079 (
  .O(mux_o_3079),
  .I0(ram16sdp_inst_502_dout[24]),
  .I1(ram16sdp_inst_510_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3080 (
  .O(mux_o_3080),
  .I0(ram16sdp_inst_518_dout[24]),
  .I1(ram16sdp_inst_526_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3081 (
  .O(mux_o_3081),
  .I0(ram16sdp_inst_534_dout[24]),
  .I1(ram16sdp_inst_542_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3082 (
  .O(mux_o_3082),
  .I0(ram16sdp_inst_550_dout[24]),
  .I1(ram16sdp_inst_558_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3083 (
  .O(mux_o_3083),
  .I0(ram16sdp_inst_566_dout[24]),
  .I1(ram16sdp_inst_574_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3084 (
  .O(mux_o_3084),
  .I0(ram16sdp_inst_582_dout[24]),
  .I1(ram16sdp_inst_590_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3085 (
  .O(mux_o_3085),
  .I0(ram16sdp_inst_598_dout[24]),
  .I1(ram16sdp_inst_606_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3086 (
  .O(mux_o_3086),
  .I0(ram16sdp_inst_614_dout[24]),
  .I1(ram16sdp_inst_622_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3087 (
  .O(mux_o_3087),
  .I0(ram16sdp_inst_630_dout[24]),
  .I1(ram16sdp_inst_638_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3088 (
  .O(mux_o_3088),
  .I0(ram16sdp_inst_646_dout[24]),
  .I1(ram16sdp_inst_654_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3089 (
  .O(mux_o_3089),
  .I0(ram16sdp_inst_662_dout[24]),
  .I1(ram16sdp_inst_670_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3090 (
  .O(mux_o_3090),
  .I0(ram16sdp_inst_678_dout[24]),
  .I1(ram16sdp_inst_686_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3091 (
  .O(mux_o_3091),
  .I0(ram16sdp_inst_694_dout[24]),
  .I1(ram16sdp_inst_702_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3092 (
  .O(mux_o_3092),
  .I0(ram16sdp_inst_710_dout[24]),
  .I1(ram16sdp_inst_718_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3093 (
  .O(mux_o_3093),
  .I0(ram16sdp_inst_726_dout[24]),
  .I1(ram16sdp_inst_734_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3094 (
  .O(mux_o_3094),
  .I0(ram16sdp_inst_742_dout[24]),
  .I1(ram16sdp_inst_750_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3095 (
  .O(mux_o_3095),
  .I0(ram16sdp_inst_758_dout[24]),
  .I1(ram16sdp_inst_766_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3096 (
  .O(mux_o_3096),
  .I0(ram16sdp_inst_774_dout[24]),
  .I1(ram16sdp_inst_782_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3097 (
  .O(mux_o_3097),
  .I0(ram16sdp_inst_790_dout[24]),
  .I1(ram16sdp_inst_798_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3098 (
  .O(mux_o_3098),
  .I0(ram16sdp_inst_806_dout[24]),
  .I1(ram16sdp_inst_814_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3099 (
  .O(mux_o_3099),
  .I0(ram16sdp_inst_822_dout[24]),
  .I1(ram16sdp_inst_830_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3100 (
  .O(mux_o_3100),
  .I0(ram16sdp_inst_838_dout[24]),
  .I1(ram16sdp_inst_846_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3101 (
  .O(mux_o_3101),
  .I0(ram16sdp_inst_854_dout[24]),
  .I1(ram16sdp_inst_862_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3102 (
  .O(mux_o_3102),
  .I0(ram16sdp_inst_870_dout[24]),
  .I1(ram16sdp_inst_878_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3103 (
  .O(mux_o_3103),
  .I0(ram16sdp_inst_886_dout[24]),
  .I1(ram16sdp_inst_894_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3104 (
  .O(mux_o_3104),
  .I0(ram16sdp_inst_902_dout[24]),
  .I1(ram16sdp_inst_910_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3105 (
  .O(mux_o_3105),
  .I0(ram16sdp_inst_918_dout[24]),
  .I1(ram16sdp_inst_926_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3106 (
  .O(mux_o_3106),
  .I0(ram16sdp_inst_934_dout[24]),
  .I1(ram16sdp_inst_942_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3107 (
  .O(mux_o_3107),
  .I0(ram16sdp_inst_950_dout[24]),
  .I1(ram16sdp_inst_958_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3108 (
  .O(mux_o_3108),
  .I0(ram16sdp_inst_966_dout[24]),
  .I1(ram16sdp_inst_974_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3109 (
  .O(mux_o_3109),
  .I0(ram16sdp_inst_982_dout[24]),
  .I1(ram16sdp_inst_990_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3110 (
  .O(mux_o_3110),
  .I0(ram16sdp_inst_998_dout[24]),
  .I1(ram16sdp_inst_1006_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3111 (
  .O(mux_o_3111),
  .I0(ram16sdp_inst_1014_dout[24]),
  .I1(ram16sdp_inst_1022_dout[24]),
  .S0(rad[4])
);
MUX2 mux_inst_3112 (
  .O(mux_o_3112),
  .I0(mux_o_3048),
  .I1(mux_o_3049),
  .S0(rad[5])
);
MUX2 mux_inst_3113 (
  .O(mux_o_3113),
  .I0(mux_o_3050),
  .I1(mux_o_3051),
  .S0(rad[5])
);
MUX2 mux_inst_3114 (
  .O(mux_o_3114),
  .I0(mux_o_3052),
  .I1(mux_o_3053),
  .S0(rad[5])
);
MUX2 mux_inst_3115 (
  .O(mux_o_3115),
  .I0(mux_o_3054),
  .I1(mux_o_3055),
  .S0(rad[5])
);
MUX2 mux_inst_3116 (
  .O(mux_o_3116),
  .I0(mux_o_3056),
  .I1(mux_o_3057),
  .S0(rad[5])
);
MUX2 mux_inst_3117 (
  .O(mux_o_3117),
  .I0(mux_o_3058),
  .I1(mux_o_3059),
  .S0(rad[5])
);
MUX2 mux_inst_3118 (
  .O(mux_o_3118),
  .I0(mux_o_3060),
  .I1(mux_o_3061),
  .S0(rad[5])
);
MUX2 mux_inst_3119 (
  .O(mux_o_3119),
  .I0(mux_o_3062),
  .I1(mux_o_3063),
  .S0(rad[5])
);
MUX2 mux_inst_3120 (
  .O(mux_o_3120),
  .I0(mux_o_3064),
  .I1(mux_o_3065),
  .S0(rad[5])
);
MUX2 mux_inst_3121 (
  .O(mux_o_3121),
  .I0(mux_o_3066),
  .I1(mux_o_3067),
  .S0(rad[5])
);
MUX2 mux_inst_3122 (
  .O(mux_o_3122),
  .I0(mux_o_3068),
  .I1(mux_o_3069),
  .S0(rad[5])
);
MUX2 mux_inst_3123 (
  .O(mux_o_3123),
  .I0(mux_o_3070),
  .I1(mux_o_3071),
  .S0(rad[5])
);
MUX2 mux_inst_3124 (
  .O(mux_o_3124),
  .I0(mux_o_3072),
  .I1(mux_o_3073),
  .S0(rad[5])
);
MUX2 mux_inst_3125 (
  .O(mux_o_3125),
  .I0(mux_o_3074),
  .I1(mux_o_3075),
  .S0(rad[5])
);
MUX2 mux_inst_3126 (
  .O(mux_o_3126),
  .I0(mux_o_3076),
  .I1(mux_o_3077),
  .S0(rad[5])
);
MUX2 mux_inst_3127 (
  .O(mux_o_3127),
  .I0(mux_o_3078),
  .I1(mux_o_3079),
  .S0(rad[5])
);
MUX2 mux_inst_3128 (
  .O(mux_o_3128),
  .I0(mux_o_3080),
  .I1(mux_o_3081),
  .S0(rad[5])
);
MUX2 mux_inst_3129 (
  .O(mux_o_3129),
  .I0(mux_o_3082),
  .I1(mux_o_3083),
  .S0(rad[5])
);
MUX2 mux_inst_3130 (
  .O(mux_o_3130),
  .I0(mux_o_3084),
  .I1(mux_o_3085),
  .S0(rad[5])
);
MUX2 mux_inst_3131 (
  .O(mux_o_3131),
  .I0(mux_o_3086),
  .I1(mux_o_3087),
  .S0(rad[5])
);
MUX2 mux_inst_3132 (
  .O(mux_o_3132),
  .I0(mux_o_3088),
  .I1(mux_o_3089),
  .S0(rad[5])
);
MUX2 mux_inst_3133 (
  .O(mux_o_3133),
  .I0(mux_o_3090),
  .I1(mux_o_3091),
  .S0(rad[5])
);
MUX2 mux_inst_3134 (
  .O(mux_o_3134),
  .I0(mux_o_3092),
  .I1(mux_o_3093),
  .S0(rad[5])
);
MUX2 mux_inst_3135 (
  .O(mux_o_3135),
  .I0(mux_o_3094),
  .I1(mux_o_3095),
  .S0(rad[5])
);
MUX2 mux_inst_3136 (
  .O(mux_o_3136),
  .I0(mux_o_3096),
  .I1(mux_o_3097),
  .S0(rad[5])
);
MUX2 mux_inst_3137 (
  .O(mux_o_3137),
  .I0(mux_o_3098),
  .I1(mux_o_3099),
  .S0(rad[5])
);
MUX2 mux_inst_3138 (
  .O(mux_o_3138),
  .I0(mux_o_3100),
  .I1(mux_o_3101),
  .S0(rad[5])
);
MUX2 mux_inst_3139 (
  .O(mux_o_3139),
  .I0(mux_o_3102),
  .I1(mux_o_3103),
  .S0(rad[5])
);
MUX2 mux_inst_3140 (
  .O(mux_o_3140),
  .I0(mux_o_3104),
  .I1(mux_o_3105),
  .S0(rad[5])
);
MUX2 mux_inst_3141 (
  .O(mux_o_3141),
  .I0(mux_o_3106),
  .I1(mux_o_3107),
  .S0(rad[5])
);
MUX2 mux_inst_3142 (
  .O(mux_o_3142),
  .I0(mux_o_3108),
  .I1(mux_o_3109),
  .S0(rad[5])
);
MUX2 mux_inst_3143 (
  .O(mux_o_3143),
  .I0(mux_o_3110),
  .I1(mux_o_3111),
  .S0(rad[5])
);
MUX2 mux_inst_3144 (
  .O(mux_o_3144),
  .I0(mux_o_3112),
  .I1(mux_o_3113),
  .S0(rad[6])
);
MUX2 mux_inst_3145 (
  .O(mux_o_3145),
  .I0(mux_o_3114),
  .I1(mux_o_3115),
  .S0(rad[6])
);
MUX2 mux_inst_3146 (
  .O(mux_o_3146),
  .I0(mux_o_3116),
  .I1(mux_o_3117),
  .S0(rad[6])
);
MUX2 mux_inst_3147 (
  .O(mux_o_3147),
  .I0(mux_o_3118),
  .I1(mux_o_3119),
  .S0(rad[6])
);
MUX2 mux_inst_3148 (
  .O(mux_o_3148),
  .I0(mux_o_3120),
  .I1(mux_o_3121),
  .S0(rad[6])
);
MUX2 mux_inst_3149 (
  .O(mux_o_3149),
  .I0(mux_o_3122),
  .I1(mux_o_3123),
  .S0(rad[6])
);
MUX2 mux_inst_3150 (
  .O(mux_o_3150),
  .I0(mux_o_3124),
  .I1(mux_o_3125),
  .S0(rad[6])
);
MUX2 mux_inst_3151 (
  .O(mux_o_3151),
  .I0(mux_o_3126),
  .I1(mux_o_3127),
  .S0(rad[6])
);
MUX2 mux_inst_3152 (
  .O(mux_o_3152),
  .I0(mux_o_3128),
  .I1(mux_o_3129),
  .S0(rad[6])
);
MUX2 mux_inst_3153 (
  .O(mux_o_3153),
  .I0(mux_o_3130),
  .I1(mux_o_3131),
  .S0(rad[6])
);
MUX2 mux_inst_3154 (
  .O(mux_o_3154),
  .I0(mux_o_3132),
  .I1(mux_o_3133),
  .S0(rad[6])
);
MUX2 mux_inst_3155 (
  .O(mux_o_3155),
  .I0(mux_o_3134),
  .I1(mux_o_3135),
  .S0(rad[6])
);
MUX2 mux_inst_3156 (
  .O(mux_o_3156),
  .I0(mux_o_3136),
  .I1(mux_o_3137),
  .S0(rad[6])
);
MUX2 mux_inst_3157 (
  .O(mux_o_3157),
  .I0(mux_o_3138),
  .I1(mux_o_3139),
  .S0(rad[6])
);
MUX2 mux_inst_3158 (
  .O(mux_o_3158),
  .I0(mux_o_3140),
  .I1(mux_o_3141),
  .S0(rad[6])
);
MUX2 mux_inst_3159 (
  .O(mux_o_3159),
  .I0(mux_o_3142),
  .I1(mux_o_3143),
  .S0(rad[6])
);
MUX2 mux_inst_3160 (
  .O(mux_o_3160),
  .I0(mux_o_3144),
  .I1(mux_o_3145),
  .S0(rad[7])
);
MUX2 mux_inst_3161 (
  .O(mux_o_3161),
  .I0(mux_o_3146),
  .I1(mux_o_3147),
  .S0(rad[7])
);
MUX2 mux_inst_3162 (
  .O(mux_o_3162),
  .I0(mux_o_3148),
  .I1(mux_o_3149),
  .S0(rad[7])
);
MUX2 mux_inst_3163 (
  .O(mux_o_3163),
  .I0(mux_o_3150),
  .I1(mux_o_3151),
  .S0(rad[7])
);
MUX2 mux_inst_3164 (
  .O(mux_o_3164),
  .I0(mux_o_3152),
  .I1(mux_o_3153),
  .S0(rad[7])
);
MUX2 mux_inst_3165 (
  .O(mux_o_3165),
  .I0(mux_o_3154),
  .I1(mux_o_3155),
  .S0(rad[7])
);
MUX2 mux_inst_3166 (
  .O(mux_o_3166),
  .I0(mux_o_3156),
  .I1(mux_o_3157),
  .S0(rad[7])
);
MUX2 mux_inst_3167 (
  .O(mux_o_3167),
  .I0(mux_o_3158),
  .I1(mux_o_3159),
  .S0(rad[7])
);
MUX2 mux_inst_3168 (
  .O(mux_o_3168),
  .I0(mux_o_3160),
  .I1(mux_o_3161),
  .S0(rad[8])
);
MUX2 mux_inst_3169 (
  .O(mux_o_3169),
  .I0(mux_o_3162),
  .I1(mux_o_3163),
  .S0(rad[8])
);
MUX2 mux_inst_3170 (
  .O(mux_o_3170),
  .I0(mux_o_3164),
  .I1(mux_o_3165),
  .S0(rad[8])
);
MUX2 mux_inst_3171 (
  .O(mux_o_3171),
  .I0(mux_o_3166),
  .I1(mux_o_3167),
  .S0(rad[8])
);
MUX2 mux_inst_3172 (
  .O(mux_o_3172),
  .I0(mux_o_3168),
  .I1(mux_o_3169),
  .S0(rad[9])
);
MUX2 mux_inst_3173 (
  .O(mux_o_3173),
  .I0(mux_o_3170),
  .I1(mux_o_3171),
  .S0(rad[9])
);
MUX2 mux_inst_3174 (
  .O(dout[24]),
  .I0(mux_o_3172),
  .I1(mux_o_3173),
  .S0(rad[10])
);
MUX2 mux_inst_3175 (
  .O(mux_o_3175),
  .I0(ram16sdp_inst_6_dout[25]),
  .I1(ram16sdp_inst_14_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3176 (
  .O(mux_o_3176),
  .I0(ram16sdp_inst_22_dout[25]),
  .I1(ram16sdp_inst_30_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3177 (
  .O(mux_o_3177),
  .I0(ram16sdp_inst_38_dout[25]),
  .I1(ram16sdp_inst_46_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3178 (
  .O(mux_o_3178),
  .I0(ram16sdp_inst_54_dout[25]),
  .I1(ram16sdp_inst_62_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3179 (
  .O(mux_o_3179),
  .I0(ram16sdp_inst_70_dout[25]),
  .I1(ram16sdp_inst_78_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3180 (
  .O(mux_o_3180),
  .I0(ram16sdp_inst_86_dout[25]),
  .I1(ram16sdp_inst_94_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3181 (
  .O(mux_o_3181),
  .I0(ram16sdp_inst_102_dout[25]),
  .I1(ram16sdp_inst_110_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3182 (
  .O(mux_o_3182),
  .I0(ram16sdp_inst_118_dout[25]),
  .I1(ram16sdp_inst_126_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3183 (
  .O(mux_o_3183),
  .I0(ram16sdp_inst_134_dout[25]),
  .I1(ram16sdp_inst_142_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3184 (
  .O(mux_o_3184),
  .I0(ram16sdp_inst_150_dout[25]),
  .I1(ram16sdp_inst_158_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3185 (
  .O(mux_o_3185),
  .I0(ram16sdp_inst_166_dout[25]),
  .I1(ram16sdp_inst_174_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3186 (
  .O(mux_o_3186),
  .I0(ram16sdp_inst_182_dout[25]),
  .I1(ram16sdp_inst_190_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3187 (
  .O(mux_o_3187),
  .I0(ram16sdp_inst_198_dout[25]),
  .I1(ram16sdp_inst_206_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3188 (
  .O(mux_o_3188),
  .I0(ram16sdp_inst_214_dout[25]),
  .I1(ram16sdp_inst_222_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3189 (
  .O(mux_o_3189),
  .I0(ram16sdp_inst_230_dout[25]),
  .I1(ram16sdp_inst_238_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3190 (
  .O(mux_o_3190),
  .I0(ram16sdp_inst_246_dout[25]),
  .I1(ram16sdp_inst_254_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3191 (
  .O(mux_o_3191),
  .I0(ram16sdp_inst_262_dout[25]),
  .I1(ram16sdp_inst_270_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3192 (
  .O(mux_o_3192),
  .I0(ram16sdp_inst_278_dout[25]),
  .I1(ram16sdp_inst_286_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3193 (
  .O(mux_o_3193),
  .I0(ram16sdp_inst_294_dout[25]),
  .I1(ram16sdp_inst_302_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3194 (
  .O(mux_o_3194),
  .I0(ram16sdp_inst_310_dout[25]),
  .I1(ram16sdp_inst_318_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3195 (
  .O(mux_o_3195),
  .I0(ram16sdp_inst_326_dout[25]),
  .I1(ram16sdp_inst_334_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3196 (
  .O(mux_o_3196),
  .I0(ram16sdp_inst_342_dout[25]),
  .I1(ram16sdp_inst_350_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3197 (
  .O(mux_o_3197),
  .I0(ram16sdp_inst_358_dout[25]),
  .I1(ram16sdp_inst_366_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3198 (
  .O(mux_o_3198),
  .I0(ram16sdp_inst_374_dout[25]),
  .I1(ram16sdp_inst_382_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3199 (
  .O(mux_o_3199),
  .I0(ram16sdp_inst_390_dout[25]),
  .I1(ram16sdp_inst_398_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3200 (
  .O(mux_o_3200),
  .I0(ram16sdp_inst_406_dout[25]),
  .I1(ram16sdp_inst_414_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3201 (
  .O(mux_o_3201),
  .I0(ram16sdp_inst_422_dout[25]),
  .I1(ram16sdp_inst_430_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3202 (
  .O(mux_o_3202),
  .I0(ram16sdp_inst_438_dout[25]),
  .I1(ram16sdp_inst_446_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3203 (
  .O(mux_o_3203),
  .I0(ram16sdp_inst_454_dout[25]),
  .I1(ram16sdp_inst_462_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3204 (
  .O(mux_o_3204),
  .I0(ram16sdp_inst_470_dout[25]),
  .I1(ram16sdp_inst_478_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3205 (
  .O(mux_o_3205),
  .I0(ram16sdp_inst_486_dout[25]),
  .I1(ram16sdp_inst_494_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3206 (
  .O(mux_o_3206),
  .I0(ram16sdp_inst_502_dout[25]),
  .I1(ram16sdp_inst_510_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3207 (
  .O(mux_o_3207),
  .I0(ram16sdp_inst_518_dout[25]),
  .I1(ram16sdp_inst_526_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3208 (
  .O(mux_o_3208),
  .I0(ram16sdp_inst_534_dout[25]),
  .I1(ram16sdp_inst_542_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3209 (
  .O(mux_o_3209),
  .I0(ram16sdp_inst_550_dout[25]),
  .I1(ram16sdp_inst_558_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3210 (
  .O(mux_o_3210),
  .I0(ram16sdp_inst_566_dout[25]),
  .I1(ram16sdp_inst_574_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3211 (
  .O(mux_o_3211),
  .I0(ram16sdp_inst_582_dout[25]),
  .I1(ram16sdp_inst_590_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3212 (
  .O(mux_o_3212),
  .I0(ram16sdp_inst_598_dout[25]),
  .I1(ram16sdp_inst_606_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3213 (
  .O(mux_o_3213),
  .I0(ram16sdp_inst_614_dout[25]),
  .I1(ram16sdp_inst_622_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3214 (
  .O(mux_o_3214),
  .I0(ram16sdp_inst_630_dout[25]),
  .I1(ram16sdp_inst_638_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3215 (
  .O(mux_o_3215),
  .I0(ram16sdp_inst_646_dout[25]),
  .I1(ram16sdp_inst_654_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3216 (
  .O(mux_o_3216),
  .I0(ram16sdp_inst_662_dout[25]),
  .I1(ram16sdp_inst_670_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3217 (
  .O(mux_o_3217),
  .I0(ram16sdp_inst_678_dout[25]),
  .I1(ram16sdp_inst_686_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3218 (
  .O(mux_o_3218),
  .I0(ram16sdp_inst_694_dout[25]),
  .I1(ram16sdp_inst_702_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3219 (
  .O(mux_o_3219),
  .I0(ram16sdp_inst_710_dout[25]),
  .I1(ram16sdp_inst_718_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3220 (
  .O(mux_o_3220),
  .I0(ram16sdp_inst_726_dout[25]),
  .I1(ram16sdp_inst_734_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3221 (
  .O(mux_o_3221),
  .I0(ram16sdp_inst_742_dout[25]),
  .I1(ram16sdp_inst_750_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3222 (
  .O(mux_o_3222),
  .I0(ram16sdp_inst_758_dout[25]),
  .I1(ram16sdp_inst_766_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3223 (
  .O(mux_o_3223),
  .I0(ram16sdp_inst_774_dout[25]),
  .I1(ram16sdp_inst_782_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3224 (
  .O(mux_o_3224),
  .I0(ram16sdp_inst_790_dout[25]),
  .I1(ram16sdp_inst_798_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3225 (
  .O(mux_o_3225),
  .I0(ram16sdp_inst_806_dout[25]),
  .I1(ram16sdp_inst_814_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3226 (
  .O(mux_o_3226),
  .I0(ram16sdp_inst_822_dout[25]),
  .I1(ram16sdp_inst_830_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3227 (
  .O(mux_o_3227),
  .I0(ram16sdp_inst_838_dout[25]),
  .I1(ram16sdp_inst_846_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3228 (
  .O(mux_o_3228),
  .I0(ram16sdp_inst_854_dout[25]),
  .I1(ram16sdp_inst_862_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3229 (
  .O(mux_o_3229),
  .I0(ram16sdp_inst_870_dout[25]),
  .I1(ram16sdp_inst_878_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3230 (
  .O(mux_o_3230),
  .I0(ram16sdp_inst_886_dout[25]),
  .I1(ram16sdp_inst_894_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3231 (
  .O(mux_o_3231),
  .I0(ram16sdp_inst_902_dout[25]),
  .I1(ram16sdp_inst_910_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3232 (
  .O(mux_o_3232),
  .I0(ram16sdp_inst_918_dout[25]),
  .I1(ram16sdp_inst_926_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3233 (
  .O(mux_o_3233),
  .I0(ram16sdp_inst_934_dout[25]),
  .I1(ram16sdp_inst_942_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3234 (
  .O(mux_o_3234),
  .I0(ram16sdp_inst_950_dout[25]),
  .I1(ram16sdp_inst_958_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3235 (
  .O(mux_o_3235),
  .I0(ram16sdp_inst_966_dout[25]),
  .I1(ram16sdp_inst_974_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3236 (
  .O(mux_o_3236),
  .I0(ram16sdp_inst_982_dout[25]),
  .I1(ram16sdp_inst_990_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3237 (
  .O(mux_o_3237),
  .I0(ram16sdp_inst_998_dout[25]),
  .I1(ram16sdp_inst_1006_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3238 (
  .O(mux_o_3238),
  .I0(ram16sdp_inst_1014_dout[25]),
  .I1(ram16sdp_inst_1022_dout[25]),
  .S0(rad[4])
);
MUX2 mux_inst_3239 (
  .O(mux_o_3239),
  .I0(mux_o_3175),
  .I1(mux_o_3176),
  .S0(rad[5])
);
MUX2 mux_inst_3240 (
  .O(mux_o_3240),
  .I0(mux_o_3177),
  .I1(mux_o_3178),
  .S0(rad[5])
);
MUX2 mux_inst_3241 (
  .O(mux_o_3241),
  .I0(mux_o_3179),
  .I1(mux_o_3180),
  .S0(rad[5])
);
MUX2 mux_inst_3242 (
  .O(mux_o_3242),
  .I0(mux_o_3181),
  .I1(mux_o_3182),
  .S0(rad[5])
);
MUX2 mux_inst_3243 (
  .O(mux_o_3243),
  .I0(mux_o_3183),
  .I1(mux_o_3184),
  .S0(rad[5])
);
MUX2 mux_inst_3244 (
  .O(mux_o_3244),
  .I0(mux_o_3185),
  .I1(mux_o_3186),
  .S0(rad[5])
);
MUX2 mux_inst_3245 (
  .O(mux_o_3245),
  .I0(mux_o_3187),
  .I1(mux_o_3188),
  .S0(rad[5])
);
MUX2 mux_inst_3246 (
  .O(mux_o_3246),
  .I0(mux_o_3189),
  .I1(mux_o_3190),
  .S0(rad[5])
);
MUX2 mux_inst_3247 (
  .O(mux_o_3247),
  .I0(mux_o_3191),
  .I1(mux_o_3192),
  .S0(rad[5])
);
MUX2 mux_inst_3248 (
  .O(mux_o_3248),
  .I0(mux_o_3193),
  .I1(mux_o_3194),
  .S0(rad[5])
);
MUX2 mux_inst_3249 (
  .O(mux_o_3249),
  .I0(mux_o_3195),
  .I1(mux_o_3196),
  .S0(rad[5])
);
MUX2 mux_inst_3250 (
  .O(mux_o_3250),
  .I0(mux_o_3197),
  .I1(mux_o_3198),
  .S0(rad[5])
);
MUX2 mux_inst_3251 (
  .O(mux_o_3251),
  .I0(mux_o_3199),
  .I1(mux_o_3200),
  .S0(rad[5])
);
MUX2 mux_inst_3252 (
  .O(mux_o_3252),
  .I0(mux_o_3201),
  .I1(mux_o_3202),
  .S0(rad[5])
);
MUX2 mux_inst_3253 (
  .O(mux_o_3253),
  .I0(mux_o_3203),
  .I1(mux_o_3204),
  .S0(rad[5])
);
MUX2 mux_inst_3254 (
  .O(mux_o_3254),
  .I0(mux_o_3205),
  .I1(mux_o_3206),
  .S0(rad[5])
);
MUX2 mux_inst_3255 (
  .O(mux_o_3255),
  .I0(mux_o_3207),
  .I1(mux_o_3208),
  .S0(rad[5])
);
MUX2 mux_inst_3256 (
  .O(mux_o_3256),
  .I0(mux_o_3209),
  .I1(mux_o_3210),
  .S0(rad[5])
);
MUX2 mux_inst_3257 (
  .O(mux_o_3257),
  .I0(mux_o_3211),
  .I1(mux_o_3212),
  .S0(rad[5])
);
MUX2 mux_inst_3258 (
  .O(mux_o_3258),
  .I0(mux_o_3213),
  .I1(mux_o_3214),
  .S0(rad[5])
);
MUX2 mux_inst_3259 (
  .O(mux_o_3259),
  .I0(mux_o_3215),
  .I1(mux_o_3216),
  .S0(rad[5])
);
MUX2 mux_inst_3260 (
  .O(mux_o_3260),
  .I0(mux_o_3217),
  .I1(mux_o_3218),
  .S0(rad[5])
);
MUX2 mux_inst_3261 (
  .O(mux_o_3261),
  .I0(mux_o_3219),
  .I1(mux_o_3220),
  .S0(rad[5])
);
MUX2 mux_inst_3262 (
  .O(mux_o_3262),
  .I0(mux_o_3221),
  .I1(mux_o_3222),
  .S0(rad[5])
);
MUX2 mux_inst_3263 (
  .O(mux_o_3263),
  .I0(mux_o_3223),
  .I1(mux_o_3224),
  .S0(rad[5])
);
MUX2 mux_inst_3264 (
  .O(mux_o_3264),
  .I0(mux_o_3225),
  .I1(mux_o_3226),
  .S0(rad[5])
);
MUX2 mux_inst_3265 (
  .O(mux_o_3265),
  .I0(mux_o_3227),
  .I1(mux_o_3228),
  .S0(rad[5])
);
MUX2 mux_inst_3266 (
  .O(mux_o_3266),
  .I0(mux_o_3229),
  .I1(mux_o_3230),
  .S0(rad[5])
);
MUX2 mux_inst_3267 (
  .O(mux_o_3267),
  .I0(mux_o_3231),
  .I1(mux_o_3232),
  .S0(rad[5])
);
MUX2 mux_inst_3268 (
  .O(mux_o_3268),
  .I0(mux_o_3233),
  .I1(mux_o_3234),
  .S0(rad[5])
);
MUX2 mux_inst_3269 (
  .O(mux_o_3269),
  .I0(mux_o_3235),
  .I1(mux_o_3236),
  .S0(rad[5])
);
MUX2 mux_inst_3270 (
  .O(mux_o_3270),
  .I0(mux_o_3237),
  .I1(mux_o_3238),
  .S0(rad[5])
);
MUX2 mux_inst_3271 (
  .O(mux_o_3271),
  .I0(mux_o_3239),
  .I1(mux_o_3240),
  .S0(rad[6])
);
MUX2 mux_inst_3272 (
  .O(mux_o_3272),
  .I0(mux_o_3241),
  .I1(mux_o_3242),
  .S0(rad[6])
);
MUX2 mux_inst_3273 (
  .O(mux_o_3273),
  .I0(mux_o_3243),
  .I1(mux_o_3244),
  .S0(rad[6])
);
MUX2 mux_inst_3274 (
  .O(mux_o_3274),
  .I0(mux_o_3245),
  .I1(mux_o_3246),
  .S0(rad[6])
);
MUX2 mux_inst_3275 (
  .O(mux_o_3275),
  .I0(mux_o_3247),
  .I1(mux_o_3248),
  .S0(rad[6])
);
MUX2 mux_inst_3276 (
  .O(mux_o_3276),
  .I0(mux_o_3249),
  .I1(mux_o_3250),
  .S0(rad[6])
);
MUX2 mux_inst_3277 (
  .O(mux_o_3277),
  .I0(mux_o_3251),
  .I1(mux_o_3252),
  .S0(rad[6])
);
MUX2 mux_inst_3278 (
  .O(mux_o_3278),
  .I0(mux_o_3253),
  .I1(mux_o_3254),
  .S0(rad[6])
);
MUX2 mux_inst_3279 (
  .O(mux_o_3279),
  .I0(mux_o_3255),
  .I1(mux_o_3256),
  .S0(rad[6])
);
MUX2 mux_inst_3280 (
  .O(mux_o_3280),
  .I0(mux_o_3257),
  .I1(mux_o_3258),
  .S0(rad[6])
);
MUX2 mux_inst_3281 (
  .O(mux_o_3281),
  .I0(mux_o_3259),
  .I1(mux_o_3260),
  .S0(rad[6])
);
MUX2 mux_inst_3282 (
  .O(mux_o_3282),
  .I0(mux_o_3261),
  .I1(mux_o_3262),
  .S0(rad[6])
);
MUX2 mux_inst_3283 (
  .O(mux_o_3283),
  .I0(mux_o_3263),
  .I1(mux_o_3264),
  .S0(rad[6])
);
MUX2 mux_inst_3284 (
  .O(mux_o_3284),
  .I0(mux_o_3265),
  .I1(mux_o_3266),
  .S0(rad[6])
);
MUX2 mux_inst_3285 (
  .O(mux_o_3285),
  .I0(mux_o_3267),
  .I1(mux_o_3268),
  .S0(rad[6])
);
MUX2 mux_inst_3286 (
  .O(mux_o_3286),
  .I0(mux_o_3269),
  .I1(mux_o_3270),
  .S0(rad[6])
);
MUX2 mux_inst_3287 (
  .O(mux_o_3287),
  .I0(mux_o_3271),
  .I1(mux_o_3272),
  .S0(rad[7])
);
MUX2 mux_inst_3288 (
  .O(mux_o_3288),
  .I0(mux_o_3273),
  .I1(mux_o_3274),
  .S0(rad[7])
);
MUX2 mux_inst_3289 (
  .O(mux_o_3289),
  .I0(mux_o_3275),
  .I1(mux_o_3276),
  .S0(rad[7])
);
MUX2 mux_inst_3290 (
  .O(mux_o_3290),
  .I0(mux_o_3277),
  .I1(mux_o_3278),
  .S0(rad[7])
);
MUX2 mux_inst_3291 (
  .O(mux_o_3291),
  .I0(mux_o_3279),
  .I1(mux_o_3280),
  .S0(rad[7])
);
MUX2 mux_inst_3292 (
  .O(mux_o_3292),
  .I0(mux_o_3281),
  .I1(mux_o_3282),
  .S0(rad[7])
);
MUX2 mux_inst_3293 (
  .O(mux_o_3293),
  .I0(mux_o_3283),
  .I1(mux_o_3284),
  .S0(rad[7])
);
MUX2 mux_inst_3294 (
  .O(mux_o_3294),
  .I0(mux_o_3285),
  .I1(mux_o_3286),
  .S0(rad[7])
);
MUX2 mux_inst_3295 (
  .O(mux_o_3295),
  .I0(mux_o_3287),
  .I1(mux_o_3288),
  .S0(rad[8])
);
MUX2 mux_inst_3296 (
  .O(mux_o_3296),
  .I0(mux_o_3289),
  .I1(mux_o_3290),
  .S0(rad[8])
);
MUX2 mux_inst_3297 (
  .O(mux_o_3297),
  .I0(mux_o_3291),
  .I1(mux_o_3292),
  .S0(rad[8])
);
MUX2 mux_inst_3298 (
  .O(mux_o_3298),
  .I0(mux_o_3293),
  .I1(mux_o_3294),
  .S0(rad[8])
);
MUX2 mux_inst_3299 (
  .O(mux_o_3299),
  .I0(mux_o_3295),
  .I1(mux_o_3296),
  .S0(rad[9])
);
MUX2 mux_inst_3300 (
  .O(mux_o_3300),
  .I0(mux_o_3297),
  .I1(mux_o_3298),
  .S0(rad[9])
);
MUX2 mux_inst_3301 (
  .O(dout[25]),
  .I0(mux_o_3299),
  .I1(mux_o_3300),
  .S0(rad[10])
);
MUX2 mux_inst_3302 (
  .O(mux_o_3302),
  .I0(ram16sdp_inst_6_dout[26]),
  .I1(ram16sdp_inst_14_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3303 (
  .O(mux_o_3303),
  .I0(ram16sdp_inst_22_dout[26]),
  .I1(ram16sdp_inst_30_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3304 (
  .O(mux_o_3304),
  .I0(ram16sdp_inst_38_dout[26]),
  .I1(ram16sdp_inst_46_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3305 (
  .O(mux_o_3305),
  .I0(ram16sdp_inst_54_dout[26]),
  .I1(ram16sdp_inst_62_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3306 (
  .O(mux_o_3306),
  .I0(ram16sdp_inst_70_dout[26]),
  .I1(ram16sdp_inst_78_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3307 (
  .O(mux_o_3307),
  .I0(ram16sdp_inst_86_dout[26]),
  .I1(ram16sdp_inst_94_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3308 (
  .O(mux_o_3308),
  .I0(ram16sdp_inst_102_dout[26]),
  .I1(ram16sdp_inst_110_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3309 (
  .O(mux_o_3309),
  .I0(ram16sdp_inst_118_dout[26]),
  .I1(ram16sdp_inst_126_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3310 (
  .O(mux_o_3310),
  .I0(ram16sdp_inst_134_dout[26]),
  .I1(ram16sdp_inst_142_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3311 (
  .O(mux_o_3311),
  .I0(ram16sdp_inst_150_dout[26]),
  .I1(ram16sdp_inst_158_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3312 (
  .O(mux_o_3312),
  .I0(ram16sdp_inst_166_dout[26]),
  .I1(ram16sdp_inst_174_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3313 (
  .O(mux_o_3313),
  .I0(ram16sdp_inst_182_dout[26]),
  .I1(ram16sdp_inst_190_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3314 (
  .O(mux_o_3314),
  .I0(ram16sdp_inst_198_dout[26]),
  .I1(ram16sdp_inst_206_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3315 (
  .O(mux_o_3315),
  .I0(ram16sdp_inst_214_dout[26]),
  .I1(ram16sdp_inst_222_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3316 (
  .O(mux_o_3316),
  .I0(ram16sdp_inst_230_dout[26]),
  .I1(ram16sdp_inst_238_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3317 (
  .O(mux_o_3317),
  .I0(ram16sdp_inst_246_dout[26]),
  .I1(ram16sdp_inst_254_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3318 (
  .O(mux_o_3318),
  .I0(ram16sdp_inst_262_dout[26]),
  .I1(ram16sdp_inst_270_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3319 (
  .O(mux_o_3319),
  .I0(ram16sdp_inst_278_dout[26]),
  .I1(ram16sdp_inst_286_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3320 (
  .O(mux_o_3320),
  .I0(ram16sdp_inst_294_dout[26]),
  .I1(ram16sdp_inst_302_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3321 (
  .O(mux_o_3321),
  .I0(ram16sdp_inst_310_dout[26]),
  .I1(ram16sdp_inst_318_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3322 (
  .O(mux_o_3322),
  .I0(ram16sdp_inst_326_dout[26]),
  .I1(ram16sdp_inst_334_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3323 (
  .O(mux_o_3323),
  .I0(ram16sdp_inst_342_dout[26]),
  .I1(ram16sdp_inst_350_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3324 (
  .O(mux_o_3324),
  .I0(ram16sdp_inst_358_dout[26]),
  .I1(ram16sdp_inst_366_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3325 (
  .O(mux_o_3325),
  .I0(ram16sdp_inst_374_dout[26]),
  .I1(ram16sdp_inst_382_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3326 (
  .O(mux_o_3326),
  .I0(ram16sdp_inst_390_dout[26]),
  .I1(ram16sdp_inst_398_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3327 (
  .O(mux_o_3327),
  .I0(ram16sdp_inst_406_dout[26]),
  .I1(ram16sdp_inst_414_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3328 (
  .O(mux_o_3328),
  .I0(ram16sdp_inst_422_dout[26]),
  .I1(ram16sdp_inst_430_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3329 (
  .O(mux_o_3329),
  .I0(ram16sdp_inst_438_dout[26]),
  .I1(ram16sdp_inst_446_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3330 (
  .O(mux_o_3330),
  .I0(ram16sdp_inst_454_dout[26]),
  .I1(ram16sdp_inst_462_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3331 (
  .O(mux_o_3331),
  .I0(ram16sdp_inst_470_dout[26]),
  .I1(ram16sdp_inst_478_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3332 (
  .O(mux_o_3332),
  .I0(ram16sdp_inst_486_dout[26]),
  .I1(ram16sdp_inst_494_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3333 (
  .O(mux_o_3333),
  .I0(ram16sdp_inst_502_dout[26]),
  .I1(ram16sdp_inst_510_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3334 (
  .O(mux_o_3334),
  .I0(ram16sdp_inst_518_dout[26]),
  .I1(ram16sdp_inst_526_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3335 (
  .O(mux_o_3335),
  .I0(ram16sdp_inst_534_dout[26]),
  .I1(ram16sdp_inst_542_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3336 (
  .O(mux_o_3336),
  .I0(ram16sdp_inst_550_dout[26]),
  .I1(ram16sdp_inst_558_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3337 (
  .O(mux_o_3337),
  .I0(ram16sdp_inst_566_dout[26]),
  .I1(ram16sdp_inst_574_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3338 (
  .O(mux_o_3338),
  .I0(ram16sdp_inst_582_dout[26]),
  .I1(ram16sdp_inst_590_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3339 (
  .O(mux_o_3339),
  .I0(ram16sdp_inst_598_dout[26]),
  .I1(ram16sdp_inst_606_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3340 (
  .O(mux_o_3340),
  .I0(ram16sdp_inst_614_dout[26]),
  .I1(ram16sdp_inst_622_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3341 (
  .O(mux_o_3341),
  .I0(ram16sdp_inst_630_dout[26]),
  .I1(ram16sdp_inst_638_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3342 (
  .O(mux_o_3342),
  .I0(ram16sdp_inst_646_dout[26]),
  .I1(ram16sdp_inst_654_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3343 (
  .O(mux_o_3343),
  .I0(ram16sdp_inst_662_dout[26]),
  .I1(ram16sdp_inst_670_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3344 (
  .O(mux_o_3344),
  .I0(ram16sdp_inst_678_dout[26]),
  .I1(ram16sdp_inst_686_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3345 (
  .O(mux_o_3345),
  .I0(ram16sdp_inst_694_dout[26]),
  .I1(ram16sdp_inst_702_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3346 (
  .O(mux_o_3346),
  .I0(ram16sdp_inst_710_dout[26]),
  .I1(ram16sdp_inst_718_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3347 (
  .O(mux_o_3347),
  .I0(ram16sdp_inst_726_dout[26]),
  .I1(ram16sdp_inst_734_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3348 (
  .O(mux_o_3348),
  .I0(ram16sdp_inst_742_dout[26]),
  .I1(ram16sdp_inst_750_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3349 (
  .O(mux_o_3349),
  .I0(ram16sdp_inst_758_dout[26]),
  .I1(ram16sdp_inst_766_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3350 (
  .O(mux_o_3350),
  .I0(ram16sdp_inst_774_dout[26]),
  .I1(ram16sdp_inst_782_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3351 (
  .O(mux_o_3351),
  .I0(ram16sdp_inst_790_dout[26]),
  .I1(ram16sdp_inst_798_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3352 (
  .O(mux_o_3352),
  .I0(ram16sdp_inst_806_dout[26]),
  .I1(ram16sdp_inst_814_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3353 (
  .O(mux_o_3353),
  .I0(ram16sdp_inst_822_dout[26]),
  .I1(ram16sdp_inst_830_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3354 (
  .O(mux_o_3354),
  .I0(ram16sdp_inst_838_dout[26]),
  .I1(ram16sdp_inst_846_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3355 (
  .O(mux_o_3355),
  .I0(ram16sdp_inst_854_dout[26]),
  .I1(ram16sdp_inst_862_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3356 (
  .O(mux_o_3356),
  .I0(ram16sdp_inst_870_dout[26]),
  .I1(ram16sdp_inst_878_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3357 (
  .O(mux_o_3357),
  .I0(ram16sdp_inst_886_dout[26]),
  .I1(ram16sdp_inst_894_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3358 (
  .O(mux_o_3358),
  .I0(ram16sdp_inst_902_dout[26]),
  .I1(ram16sdp_inst_910_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3359 (
  .O(mux_o_3359),
  .I0(ram16sdp_inst_918_dout[26]),
  .I1(ram16sdp_inst_926_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3360 (
  .O(mux_o_3360),
  .I0(ram16sdp_inst_934_dout[26]),
  .I1(ram16sdp_inst_942_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3361 (
  .O(mux_o_3361),
  .I0(ram16sdp_inst_950_dout[26]),
  .I1(ram16sdp_inst_958_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3362 (
  .O(mux_o_3362),
  .I0(ram16sdp_inst_966_dout[26]),
  .I1(ram16sdp_inst_974_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3363 (
  .O(mux_o_3363),
  .I0(ram16sdp_inst_982_dout[26]),
  .I1(ram16sdp_inst_990_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3364 (
  .O(mux_o_3364),
  .I0(ram16sdp_inst_998_dout[26]),
  .I1(ram16sdp_inst_1006_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3365 (
  .O(mux_o_3365),
  .I0(ram16sdp_inst_1014_dout[26]),
  .I1(ram16sdp_inst_1022_dout[26]),
  .S0(rad[4])
);
MUX2 mux_inst_3366 (
  .O(mux_o_3366),
  .I0(mux_o_3302),
  .I1(mux_o_3303),
  .S0(rad[5])
);
MUX2 mux_inst_3367 (
  .O(mux_o_3367),
  .I0(mux_o_3304),
  .I1(mux_o_3305),
  .S0(rad[5])
);
MUX2 mux_inst_3368 (
  .O(mux_o_3368),
  .I0(mux_o_3306),
  .I1(mux_o_3307),
  .S0(rad[5])
);
MUX2 mux_inst_3369 (
  .O(mux_o_3369),
  .I0(mux_o_3308),
  .I1(mux_o_3309),
  .S0(rad[5])
);
MUX2 mux_inst_3370 (
  .O(mux_o_3370),
  .I0(mux_o_3310),
  .I1(mux_o_3311),
  .S0(rad[5])
);
MUX2 mux_inst_3371 (
  .O(mux_o_3371),
  .I0(mux_o_3312),
  .I1(mux_o_3313),
  .S0(rad[5])
);
MUX2 mux_inst_3372 (
  .O(mux_o_3372),
  .I0(mux_o_3314),
  .I1(mux_o_3315),
  .S0(rad[5])
);
MUX2 mux_inst_3373 (
  .O(mux_o_3373),
  .I0(mux_o_3316),
  .I1(mux_o_3317),
  .S0(rad[5])
);
MUX2 mux_inst_3374 (
  .O(mux_o_3374),
  .I0(mux_o_3318),
  .I1(mux_o_3319),
  .S0(rad[5])
);
MUX2 mux_inst_3375 (
  .O(mux_o_3375),
  .I0(mux_o_3320),
  .I1(mux_o_3321),
  .S0(rad[5])
);
MUX2 mux_inst_3376 (
  .O(mux_o_3376),
  .I0(mux_o_3322),
  .I1(mux_o_3323),
  .S0(rad[5])
);
MUX2 mux_inst_3377 (
  .O(mux_o_3377),
  .I0(mux_o_3324),
  .I1(mux_o_3325),
  .S0(rad[5])
);
MUX2 mux_inst_3378 (
  .O(mux_o_3378),
  .I0(mux_o_3326),
  .I1(mux_o_3327),
  .S0(rad[5])
);
MUX2 mux_inst_3379 (
  .O(mux_o_3379),
  .I0(mux_o_3328),
  .I1(mux_o_3329),
  .S0(rad[5])
);
MUX2 mux_inst_3380 (
  .O(mux_o_3380),
  .I0(mux_o_3330),
  .I1(mux_o_3331),
  .S0(rad[5])
);
MUX2 mux_inst_3381 (
  .O(mux_o_3381),
  .I0(mux_o_3332),
  .I1(mux_o_3333),
  .S0(rad[5])
);
MUX2 mux_inst_3382 (
  .O(mux_o_3382),
  .I0(mux_o_3334),
  .I1(mux_o_3335),
  .S0(rad[5])
);
MUX2 mux_inst_3383 (
  .O(mux_o_3383),
  .I0(mux_o_3336),
  .I1(mux_o_3337),
  .S0(rad[5])
);
MUX2 mux_inst_3384 (
  .O(mux_o_3384),
  .I0(mux_o_3338),
  .I1(mux_o_3339),
  .S0(rad[5])
);
MUX2 mux_inst_3385 (
  .O(mux_o_3385),
  .I0(mux_o_3340),
  .I1(mux_o_3341),
  .S0(rad[5])
);
MUX2 mux_inst_3386 (
  .O(mux_o_3386),
  .I0(mux_o_3342),
  .I1(mux_o_3343),
  .S0(rad[5])
);
MUX2 mux_inst_3387 (
  .O(mux_o_3387),
  .I0(mux_o_3344),
  .I1(mux_o_3345),
  .S0(rad[5])
);
MUX2 mux_inst_3388 (
  .O(mux_o_3388),
  .I0(mux_o_3346),
  .I1(mux_o_3347),
  .S0(rad[5])
);
MUX2 mux_inst_3389 (
  .O(mux_o_3389),
  .I0(mux_o_3348),
  .I1(mux_o_3349),
  .S0(rad[5])
);
MUX2 mux_inst_3390 (
  .O(mux_o_3390),
  .I0(mux_o_3350),
  .I1(mux_o_3351),
  .S0(rad[5])
);
MUX2 mux_inst_3391 (
  .O(mux_o_3391),
  .I0(mux_o_3352),
  .I1(mux_o_3353),
  .S0(rad[5])
);
MUX2 mux_inst_3392 (
  .O(mux_o_3392),
  .I0(mux_o_3354),
  .I1(mux_o_3355),
  .S0(rad[5])
);
MUX2 mux_inst_3393 (
  .O(mux_o_3393),
  .I0(mux_o_3356),
  .I1(mux_o_3357),
  .S0(rad[5])
);
MUX2 mux_inst_3394 (
  .O(mux_o_3394),
  .I0(mux_o_3358),
  .I1(mux_o_3359),
  .S0(rad[5])
);
MUX2 mux_inst_3395 (
  .O(mux_o_3395),
  .I0(mux_o_3360),
  .I1(mux_o_3361),
  .S0(rad[5])
);
MUX2 mux_inst_3396 (
  .O(mux_o_3396),
  .I0(mux_o_3362),
  .I1(mux_o_3363),
  .S0(rad[5])
);
MUX2 mux_inst_3397 (
  .O(mux_o_3397),
  .I0(mux_o_3364),
  .I1(mux_o_3365),
  .S0(rad[5])
);
MUX2 mux_inst_3398 (
  .O(mux_o_3398),
  .I0(mux_o_3366),
  .I1(mux_o_3367),
  .S0(rad[6])
);
MUX2 mux_inst_3399 (
  .O(mux_o_3399),
  .I0(mux_o_3368),
  .I1(mux_o_3369),
  .S0(rad[6])
);
MUX2 mux_inst_3400 (
  .O(mux_o_3400),
  .I0(mux_o_3370),
  .I1(mux_o_3371),
  .S0(rad[6])
);
MUX2 mux_inst_3401 (
  .O(mux_o_3401),
  .I0(mux_o_3372),
  .I1(mux_o_3373),
  .S0(rad[6])
);
MUX2 mux_inst_3402 (
  .O(mux_o_3402),
  .I0(mux_o_3374),
  .I1(mux_o_3375),
  .S0(rad[6])
);
MUX2 mux_inst_3403 (
  .O(mux_o_3403),
  .I0(mux_o_3376),
  .I1(mux_o_3377),
  .S0(rad[6])
);
MUX2 mux_inst_3404 (
  .O(mux_o_3404),
  .I0(mux_o_3378),
  .I1(mux_o_3379),
  .S0(rad[6])
);
MUX2 mux_inst_3405 (
  .O(mux_o_3405),
  .I0(mux_o_3380),
  .I1(mux_o_3381),
  .S0(rad[6])
);
MUX2 mux_inst_3406 (
  .O(mux_o_3406),
  .I0(mux_o_3382),
  .I1(mux_o_3383),
  .S0(rad[6])
);
MUX2 mux_inst_3407 (
  .O(mux_o_3407),
  .I0(mux_o_3384),
  .I1(mux_o_3385),
  .S0(rad[6])
);
MUX2 mux_inst_3408 (
  .O(mux_o_3408),
  .I0(mux_o_3386),
  .I1(mux_o_3387),
  .S0(rad[6])
);
MUX2 mux_inst_3409 (
  .O(mux_o_3409),
  .I0(mux_o_3388),
  .I1(mux_o_3389),
  .S0(rad[6])
);
MUX2 mux_inst_3410 (
  .O(mux_o_3410),
  .I0(mux_o_3390),
  .I1(mux_o_3391),
  .S0(rad[6])
);
MUX2 mux_inst_3411 (
  .O(mux_o_3411),
  .I0(mux_o_3392),
  .I1(mux_o_3393),
  .S0(rad[6])
);
MUX2 mux_inst_3412 (
  .O(mux_o_3412),
  .I0(mux_o_3394),
  .I1(mux_o_3395),
  .S0(rad[6])
);
MUX2 mux_inst_3413 (
  .O(mux_o_3413),
  .I0(mux_o_3396),
  .I1(mux_o_3397),
  .S0(rad[6])
);
MUX2 mux_inst_3414 (
  .O(mux_o_3414),
  .I0(mux_o_3398),
  .I1(mux_o_3399),
  .S0(rad[7])
);
MUX2 mux_inst_3415 (
  .O(mux_o_3415),
  .I0(mux_o_3400),
  .I1(mux_o_3401),
  .S0(rad[7])
);
MUX2 mux_inst_3416 (
  .O(mux_o_3416),
  .I0(mux_o_3402),
  .I1(mux_o_3403),
  .S0(rad[7])
);
MUX2 mux_inst_3417 (
  .O(mux_o_3417),
  .I0(mux_o_3404),
  .I1(mux_o_3405),
  .S0(rad[7])
);
MUX2 mux_inst_3418 (
  .O(mux_o_3418),
  .I0(mux_o_3406),
  .I1(mux_o_3407),
  .S0(rad[7])
);
MUX2 mux_inst_3419 (
  .O(mux_o_3419),
  .I0(mux_o_3408),
  .I1(mux_o_3409),
  .S0(rad[7])
);
MUX2 mux_inst_3420 (
  .O(mux_o_3420),
  .I0(mux_o_3410),
  .I1(mux_o_3411),
  .S0(rad[7])
);
MUX2 mux_inst_3421 (
  .O(mux_o_3421),
  .I0(mux_o_3412),
  .I1(mux_o_3413),
  .S0(rad[7])
);
MUX2 mux_inst_3422 (
  .O(mux_o_3422),
  .I0(mux_o_3414),
  .I1(mux_o_3415),
  .S0(rad[8])
);
MUX2 mux_inst_3423 (
  .O(mux_o_3423),
  .I0(mux_o_3416),
  .I1(mux_o_3417),
  .S0(rad[8])
);
MUX2 mux_inst_3424 (
  .O(mux_o_3424),
  .I0(mux_o_3418),
  .I1(mux_o_3419),
  .S0(rad[8])
);
MUX2 mux_inst_3425 (
  .O(mux_o_3425),
  .I0(mux_o_3420),
  .I1(mux_o_3421),
  .S0(rad[8])
);
MUX2 mux_inst_3426 (
  .O(mux_o_3426),
  .I0(mux_o_3422),
  .I1(mux_o_3423),
  .S0(rad[9])
);
MUX2 mux_inst_3427 (
  .O(mux_o_3427),
  .I0(mux_o_3424),
  .I1(mux_o_3425),
  .S0(rad[9])
);
MUX2 mux_inst_3428 (
  .O(dout[26]),
  .I0(mux_o_3426),
  .I1(mux_o_3427),
  .S0(rad[10])
);
MUX2 mux_inst_3429 (
  .O(mux_o_3429),
  .I0(ram16sdp_inst_6_dout[27]),
  .I1(ram16sdp_inst_14_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3430 (
  .O(mux_o_3430),
  .I0(ram16sdp_inst_22_dout[27]),
  .I1(ram16sdp_inst_30_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3431 (
  .O(mux_o_3431),
  .I0(ram16sdp_inst_38_dout[27]),
  .I1(ram16sdp_inst_46_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3432 (
  .O(mux_o_3432),
  .I0(ram16sdp_inst_54_dout[27]),
  .I1(ram16sdp_inst_62_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3433 (
  .O(mux_o_3433),
  .I0(ram16sdp_inst_70_dout[27]),
  .I1(ram16sdp_inst_78_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3434 (
  .O(mux_o_3434),
  .I0(ram16sdp_inst_86_dout[27]),
  .I1(ram16sdp_inst_94_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3435 (
  .O(mux_o_3435),
  .I0(ram16sdp_inst_102_dout[27]),
  .I1(ram16sdp_inst_110_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3436 (
  .O(mux_o_3436),
  .I0(ram16sdp_inst_118_dout[27]),
  .I1(ram16sdp_inst_126_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3437 (
  .O(mux_o_3437),
  .I0(ram16sdp_inst_134_dout[27]),
  .I1(ram16sdp_inst_142_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3438 (
  .O(mux_o_3438),
  .I0(ram16sdp_inst_150_dout[27]),
  .I1(ram16sdp_inst_158_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3439 (
  .O(mux_o_3439),
  .I0(ram16sdp_inst_166_dout[27]),
  .I1(ram16sdp_inst_174_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3440 (
  .O(mux_o_3440),
  .I0(ram16sdp_inst_182_dout[27]),
  .I1(ram16sdp_inst_190_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3441 (
  .O(mux_o_3441),
  .I0(ram16sdp_inst_198_dout[27]),
  .I1(ram16sdp_inst_206_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3442 (
  .O(mux_o_3442),
  .I0(ram16sdp_inst_214_dout[27]),
  .I1(ram16sdp_inst_222_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3443 (
  .O(mux_o_3443),
  .I0(ram16sdp_inst_230_dout[27]),
  .I1(ram16sdp_inst_238_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3444 (
  .O(mux_o_3444),
  .I0(ram16sdp_inst_246_dout[27]),
  .I1(ram16sdp_inst_254_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3445 (
  .O(mux_o_3445),
  .I0(ram16sdp_inst_262_dout[27]),
  .I1(ram16sdp_inst_270_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3446 (
  .O(mux_o_3446),
  .I0(ram16sdp_inst_278_dout[27]),
  .I1(ram16sdp_inst_286_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3447 (
  .O(mux_o_3447),
  .I0(ram16sdp_inst_294_dout[27]),
  .I1(ram16sdp_inst_302_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3448 (
  .O(mux_o_3448),
  .I0(ram16sdp_inst_310_dout[27]),
  .I1(ram16sdp_inst_318_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3449 (
  .O(mux_o_3449),
  .I0(ram16sdp_inst_326_dout[27]),
  .I1(ram16sdp_inst_334_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3450 (
  .O(mux_o_3450),
  .I0(ram16sdp_inst_342_dout[27]),
  .I1(ram16sdp_inst_350_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3451 (
  .O(mux_o_3451),
  .I0(ram16sdp_inst_358_dout[27]),
  .I1(ram16sdp_inst_366_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3452 (
  .O(mux_o_3452),
  .I0(ram16sdp_inst_374_dout[27]),
  .I1(ram16sdp_inst_382_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3453 (
  .O(mux_o_3453),
  .I0(ram16sdp_inst_390_dout[27]),
  .I1(ram16sdp_inst_398_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3454 (
  .O(mux_o_3454),
  .I0(ram16sdp_inst_406_dout[27]),
  .I1(ram16sdp_inst_414_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3455 (
  .O(mux_o_3455),
  .I0(ram16sdp_inst_422_dout[27]),
  .I1(ram16sdp_inst_430_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3456 (
  .O(mux_o_3456),
  .I0(ram16sdp_inst_438_dout[27]),
  .I1(ram16sdp_inst_446_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3457 (
  .O(mux_o_3457),
  .I0(ram16sdp_inst_454_dout[27]),
  .I1(ram16sdp_inst_462_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3458 (
  .O(mux_o_3458),
  .I0(ram16sdp_inst_470_dout[27]),
  .I1(ram16sdp_inst_478_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3459 (
  .O(mux_o_3459),
  .I0(ram16sdp_inst_486_dout[27]),
  .I1(ram16sdp_inst_494_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3460 (
  .O(mux_o_3460),
  .I0(ram16sdp_inst_502_dout[27]),
  .I1(ram16sdp_inst_510_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3461 (
  .O(mux_o_3461),
  .I0(ram16sdp_inst_518_dout[27]),
  .I1(ram16sdp_inst_526_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3462 (
  .O(mux_o_3462),
  .I0(ram16sdp_inst_534_dout[27]),
  .I1(ram16sdp_inst_542_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3463 (
  .O(mux_o_3463),
  .I0(ram16sdp_inst_550_dout[27]),
  .I1(ram16sdp_inst_558_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3464 (
  .O(mux_o_3464),
  .I0(ram16sdp_inst_566_dout[27]),
  .I1(ram16sdp_inst_574_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3465 (
  .O(mux_o_3465),
  .I0(ram16sdp_inst_582_dout[27]),
  .I1(ram16sdp_inst_590_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3466 (
  .O(mux_o_3466),
  .I0(ram16sdp_inst_598_dout[27]),
  .I1(ram16sdp_inst_606_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3467 (
  .O(mux_o_3467),
  .I0(ram16sdp_inst_614_dout[27]),
  .I1(ram16sdp_inst_622_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3468 (
  .O(mux_o_3468),
  .I0(ram16sdp_inst_630_dout[27]),
  .I1(ram16sdp_inst_638_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3469 (
  .O(mux_o_3469),
  .I0(ram16sdp_inst_646_dout[27]),
  .I1(ram16sdp_inst_654_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3470 (
  .O(mux_o_3470),
  .I0(ram16sdp_inst_662_dout[27]),
  .I1(ram16sdp_inst_670_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3471 (
  .O(mux_o_3471),
  .I0(ram16sdp_inst_678_dout[27]),
  .I1(ram16sdp_inst_686_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3472 (
  .O(mux_o_3472),
  .I0(ram16sdp_inst_694_dout[27]),
  .I1(ram16sdp_inst_702_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3473 (
  .O(mux_o_3473),
  .I0(ram16sdp_inst_710_dout[27]),
  .I1(ram16sdp_inst_718_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3474 (
  .O(mux_o_3474),
  .I0(ram16sdp_inst_726_dout[27]),
  .I1(ram16sdp_inst_734_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3475 (
  .O(mux_o_3475),
  .I0(ram16sdp_inst_742_dout[27]),
  .I1(ram16sdp_inst_750_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3476 (
  .O(mux_o_3476),
  .I0(ram16sdp_inst_758_dout[27]),
  .I1(ram16sdp_inst_766_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3477 (
  .O(mux_o_3477),
  .I0(ram16sdp_inst_774_dout[27]),
  .I1(ram16sdp_inst_782_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3478 (
  .O(mux_o_3478),
  .I0(ram16sdp_inst_790_dout[27]),
  .I1(ram16sdp_inst_798_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3479 (
  .O(mux_o_3479),
  .I0(ram16sdp_inst_806_dout[27]),
  .I1(ram16sdp_inst_814_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3480 (
  .O(mux_o_3480),
  .I0(ram16sdp_inst_822_dout[27]),
  .I1(ram16sdp_inst_830_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3481 (
  .O(mux_o_3481),
  .I0(ram16sdp_inst_838_dout[27]),
  .I1(ram16sdp_inst_846_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3482 (
  .O(mux_o_3482),
  .I0(ram16sdp_inst_854_dout[27]),
  .I1(ram16sdp_inst_862_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3483 (
  .O(mux_o_3483),
  .I0(ram16sdp_inst_870_dout[27]),
  .I1(ram16sdp_inst_878_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3484 (
  .O(mux_o_3484),
  .I0(ram16sdp_inst_886_dout[27]),
  .I1(ram16sdp_inst_894_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3485 (
  .O(mux_o_3485),
  .I0(ram16sdp_inst_902_dout[27]),
  .I1(ram16sdp_inst_910_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3486 (
  .O(mux_o_3486),
  .I0(ram16sdp_inst_918_dout[27]),
  .I1(ram16sdp_inst_926_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3487 (
  .O(mux_o_3487),
  .I0(ram16sdp_inst_934_dout[27]),
  .I1(ram16sdp_inst_942_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3488 (
  .O(mux_o_3488),
  .I0(ram16sdp_inst_950_dout[27]),
  .I1(ram16sdp_inst_958_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3489 (
  .O(mux_o_3489),
  .I0(ram16sdp_inst_966_dout[27]),
  .I1(ram16sdp_inst_974_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3490 (
  .O(mux_o_3490),
  .I0(ram16sdp_inst_982_dout[27]),
  .I1(ram16sdp_inst_990_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3491 (
  .O(mux_o_3491),
  .I0(ram16sdp_inst_998_dout[27]),
  .I1(ram16sdp_inst_1006_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3492 (
  .O(mux_o_3492),
  .I0(ram16sdp_inst_1014_dout[27]),
  .I1(ram16sdp_inst_1022_dout[27]),
  .S0(rad[4])
);
MUX2 mux_inst_3493 (
  .O(mux_o_3493),
  .I0(mux_o_3429),
  .I1(mux_o_3430),
  .S0(rad[5])
);
MUX2 mux_inst_3494 (
  .O(mux_o_3494),
  .I0(mux_o_3431),
  .I1(mux_o_3432),
  .S0(rad[5])
);
MUX2 mux_inst_3495 (
  .O(mux_o_3495),
  .I0(mux_o_3433),
  .I1(mux_o_3434),
  .S0(rad[5])
);
MUX2 mux_inst_3496 (
  .O(mux_o_3496),
  .I0(mux_o_3435),
  .I1(mux_o_3436),
  .S0(rad[5])
);
MUX2 mux_inst_3497 (
  .O(mux_o_3497),
  .I0(mux_o_3437),
  .I1(mux_o_3438),
  .S0(rad[5])
);
MUX2 mux_inst_3498 (
  .O(mux_o_3498),
  .I0(mux_o_3439),
  .I1(mux_o_3440),
  .S0(rad[5])
);
MUX2 mux_inst_3499 (
  .O(mux_o_3499),
  .I0(mux_o_3441),
  .I1(mux_o_3442),
  .S0(rad[5])
);
MUX2 mux_inst_3500 (
  .O(mux_o_3500),
  .I0(mux_o_3443),
  .I1(mux_o_3444),
  .S0(rad[5])
);
MUX2 mux_inst_3501 (
  .O(mux_o_3501),
  .I0(mux_o_3445),
  .I1(mux_o_3446),
  .S0(rad[5])
);
MUX2 mux_inst_3502 (
  .O(mux_o_3502),
  .I0(mux_o_3447),
  .I1(mux_o_3448),
  .S0(rad[5])
);
MUX2 mux_inst_3503 (
  .O(mux_o_3503),
  .I0(mux_o_3449),
  .I1(mux_o_3450),
  .S0(rad[5])
);
MUX2 mux_inst_3504 (
  .O(mux_o_3504),
  .I0(mux_o_3451),
  .I1(mux_o_3452),
  .S0(rad[5])
);
MUX2 mux_inst_3505 (
  .O(mux_o_3505),
  .I0(mux_o_3453),
  .I1(mux_o_3454),
  .S0(rad[5])
);
MUX2 mux_inst_3506 (
  .O(mux_o_3506),
  .I0(mux_o_3455),
  .I1(mux_o_3456),
  .S0(rad[5])
);
MUX2 mux_inst_3507 (
  .O(mux_o_3507),
  .I0(mux_o_3457),
  .I1(mux_o_3458),
  .S0(rad[5])
);
MUX2 mux_inst_3508 (
  .O(mux_o_3508),
  .I0(mux_o_3459),
  .I1(mux_o_3460),
  .S0(rad[5])
);
MUX2 mux_inst_3509 (
  .O(mux_o_3509),
  .I0(mux_o_3461),
  .I1(mux_o_3462),
  .S0(rad[5])
);
MUX2 mux_inst_3510 (
  .O(mux_o_3510),
  .I0(mux_o_3463),
  .I1(mux_o_3464),
  .S0(rad[5])
);
MUX2 mux_inst_3511 (
  .O(mux_o_3511),
  .I0(mux_o_3465),
  .I1(mux_o_3466),
  .S0(rad[5])
);
MUX2 mux_inst_3512 (
  .O(mux_o_3512),
  .I0(mux_o_3467),
  .I1(mux_o_3468),
  .S0(rad[5])
);
MUX2 mux_inst_3513 (
  .O(mux_o_3513),
  .I0(mux_o_3469),
  .I1(mux_o_3470),
  .S0(rad[5])
);
MUX2 mux_inst_3514 (
  .O(mux_o_3514),
  .I0(mux_o_3471),
  .I1(mux_o_3472),
  .S0(rad[5])
);
MUX2 mux_inst_3515 (
  .O(mux_o_3515),
  .I0(mux_o_3473),
  .I1(mux_o_3474),
  .S0(rad[5])
);
MUX2 mux_inst_3516 (
  .O(mux_o_3516),
  .I0(mux_o_3475),
  .I1(mux_o_3476),
  .S0(rad[5])
);
MUX2 mux_inst_3517 (
  .O(mux_o_3517),
  .I0(mux_o_3477),
  .I1(mux_o_3478),
  .S0(rad[5])
);
MUX2 mux_inst_3518 (
  .O(mux_o_3518),
  .I0(mux_o_3479),
  .I1(mux_o_3480),
  .S0(rad[5])
);
MUX2 mux_inst_3519 (
  .O(mux_o_3519),
  .I0(mux_o_3481),
  .I1(mux_o_3482),
  .S0(rad[5])
);
MUX2 mux_inst_3520 (
  .O(mux_o_3520),
  .I0(mux_o_3483),
  .I1(mux_o_3484),
  .S0(rad[5])
);
MUX2 mux_inst_3521 (
  .O(mux_o_3521),
  .I0(mux_o_3485),
  .I1(mux_o_3486),
  .S0(rad[5])
);
MUX2 mux_inst_3522 (
  .O(mux_o_3522),
  .I0(mux_o_3487),
  .I1(mux_o_3488),
  .S0(rad[5])
);
MUX2 mux_inst_3523 (
  .O(mux_o_3523),
  .I0(mux_o_3489),
  .I1(mux_o_3490),
  .S0(rad[5])
);
MUX2 mux_inst_3524 (
  .O(mux_o_3524),
  .I0(mux_o_3491),
  .I1(mux_o_3492),
  .S0(rad[5])
);
MUX2 mux_inst_3525 (
  .O(mux_o_3525),
  .I0(mux_o_3493),
  .I1(mux_o_3494),
  .S0(rad[6])
);
MUX2 mux_inst_3526 (
  .O(mux_o_3526),
  .I0(mux_o_3495),
  .I1(mux_o_3496),
  .S0(rad[6])
);
MUX2 mux_inst_3527 (
  .O(mux_o_3527),
  .I0(mux_o_3497),
  .I1(mux_o_3498),
  .S0(rad[6])
);
MUX2 mux_inst_3528 (
  .O(mux_o_3528),
  .I0(mux_o_3499),
  .I1(mux_o_3500),
  .S0(rad[6])
);
MUX2 mux_inst_3529 (
  .O(mux_o_3529),
  .I0(mux_o_3501),
  .I1(mux_o_3502),
  .S0(rad[6])
);
MUX2 mux_inst_3530 (
  .O(mux_o_3530),
  .I0(mux_o_3503),
  .I1(mux_o_3504),
  .S0(rad[6])
);
MUX2 mux_inst_3531 (
  .O(mux_o_3531),
  .I0(mux_o_3505),
  .I1(mux_o_3506),
  .S0(rad[6])
);
MUX2 mux_inst_3532 (
  .O(mux_o_3532),
  .I0(mux_o_3507),
  .I1(mux_o_3508),
  .S0(rad[6])
);
MUX2 mux_inst_3533 (
  .O(mux_o_3533),
  .I0(mux_o_3509),
  .I1(mux_o_3510),
  .S0(rad[6])
);
MUX2 mux_inst_3534 (
  .O(mux_o_3534),
  .I0(mux_o_3511),
  .I1(mux_o_3512),
  .S0(rad[6])
);
MUX2 mux_inst_3535 (
  .O(mux_o_3535),
  .I0(mux_o_3513),
  .I1(mux_o_3514),
  .S0(rad[6])
);
MUX2 mux_inst_3536 (
  .O(mux_o_3536),
  .I0(mux_o_3515),
  .I1(mux_o_3516),
  .S0(rad[6])
);
MUX2 mux_inst_3537 (
  .O(mux_o_3537),
  .I0(mux_o_3517),
  .I1(mux_o_3518),
  .S0(rad[6])
);
MUX2 mux_inst_3538 (
  .O(mux_o_3538),
  .I0(mux_o_3519),
  .I1(mux_o_3520),
  .S0(rad[6])
);
MUX2 mux_inst_3539 (
  .O(mux_o_3539),
  .I0(mux_o_3521),
  .I1(mux_o_3522),
  .S0(rad[6])
);
MUX2 mux_inst_3540 (
  .O(mux_o_3540),
  .I0(mux_o_3523),
  .I1(mux_o_3524),
  .S0(rad[6])
);
MUX2 mux_inst_3541 (
  .O(mux_o_3541),
  .I0(mux_o_3525),
  .I1(mux_o_3526),
  .S0(rad[7])
);
MUX2 mux_inst_3542 (
  .O(mux_o_3542),
  .I0(mux_o_3527),
  .I1(mux_o_3528),
  .S0(rad[7])
);
MUX2 mux_inst_3543 (
  .O(mux_o_3543),
  .I0(mux_o_3529),
  .I1(mux_o_3530),
  .S0(rad[7])
);
MUX2 mux_inst_3544 (
  .O(mux_o_3544),
  .I0(mux_o_3531),
  .I1(mux_o_3532),
  .S0(rad[7])
);
MUX2 mux_inst_3545 (
  .O(mux_o_3545),
  .I0(mux_o_3533),
  .I1(mux_o_3534),
  .S0(rad[7])
);
MUX2 mux_inst_3546 (
  .O(mux_o_3546),
  .I0(mux_o_3535),
  .I1(mux_o_3536),
  .S0(rad[7])
);
MUX2 mux_inst_3547 (
  .O(mux_o_3547),
  .I0(mux_o_3537),
  .I1(mux_o_3538),
  .S0(rad[7])
);
MUX2 mux_inst_3548 (
  .O(mux_o_3548),
  .I0(mux_o_3539),
  .I1(mux_o_3540),
  .S0(rad[7])
);
MUX2 mux_inst_3549 (
  .O(mux_o_3549),
  .I0(mux_o_3541),
  .I1(mux_o_3542),
  .S0(rad[8])
);
MUX2 mux_inst_3550 (
  .O(mux_o_3550),
  .I0(mux_o_3543),
  .I1(mux_o_3544),
  .S0(rad[8])
);
MUX2 mux_inst_3551 (
  .O(mux_o_3551),
  .I0(mux_o_3545),
  .I1(mux_o_3546),
  .S0(rad[8])
);
MUX2 mux_inst_3552 (
  .O(mux_o_3552),
  .I0(mux_o_3547),
  .I1(mux_o_3548),
  .S0(rad[8])
);
MUX2 mux_inst_3553 (
  .O(mux_o_3553),
  .I0(mux_o_3549),
  .I1(mux_o_3550),
  .S0(rad[9])
);
MUX2 mux_inst_3554 (
  .O(mux_o_3554),
  .I0(mux_o_3551),
  .I1(mux_o_3552),
  .S0(rad[9])
);
MUX2 mux_inst_3555 (
  .O(dout[27]),
  .I0(mux_o_3553),
  .I1(mux_o_3554),
  .S0(rad[10])
);
MUX2 mux_inst_3556 (
  .O(mux_o_3556),
  .I0(ram16sdp_inst_7_dout[28]),
  .I1(ram16sdp_inst_15_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3557 (
  .O(mux_o_3557),
  .I0(ram16sdp_inst_23_dout[28]),
  .I1(ram16sdp_inst_31_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3558 (
  .O(mux_o_3558),
  .I0(ram16sdp_inst_39_dout[28]),
  .I1(ram16sdp_inst_47_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3559 (
  .O(mux_o_3559),
  .I0(ram16sdp_inst_55_dout[28]),
  .I1(ram16sdp_inst_63_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3560 (
  .O(mux_o_3560),
  .I0(ram16sdp_inst_71_dout[28]),
  .I1(ram16sdp_inst_79_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3561 (
  .O(mux_o_3561),
  .I0(ram16sdp_inst_87_dout[28]),
  .I1(ram16sdp_inst_95_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3562 (
  .O(mux_o_3562),
  .I0(ram16sdp_inst_103_dout[28]),
  .I1(ram16sdp_inst_111_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3563 (
  .O(mux_o_3563),
  .I0(ram16sdp_inst_119_dout[28]),
  .I1(ram16sdp_inst_127_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3564 (
  .O(mux_o_3564),
  .I0(ram16sdp_inst_135_dout[28]),
  .I1(ram16sdp_inst_143_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3565 (
  .O(mux_o_3565),
  .I0(ram16sdp_inst_151_dout[28]),
  .I1(ram16sdp_inst_159_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3566 (
  .O(mux_o_3566),
  .I0(ram16sdp_inst_167_dout[28]),
  .I1(ram16sdp_inst_175_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3567 (
  .O(mux_o_3567),
  .I0(ram16sdp_inst_183_dout[28]),
  .I1(ram16sdp_inst_191_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3568 (
  .O(mux_o_3568),
  .I0(ram16sdp_inst_199_dout[28]),
  .I1(ram16sdp_inst_207_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3569 (
  .O(mux_o_3569),
  .I0(ram16sdp_inst_215_dout[28]),
  .I1(ram16sdp_inst_223_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3570 (
  .O(mux_o_3570),
  .I0(ram16sdp_inst_231_dout[28]),
  .I1(ram16sdp_inst_239_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3571 (
  .O(mux_o_3571),
  .I0(ram16sdp_inst_247_dout[28]),
  .I1(ram16sdp_inst_255_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3572 (
  .O(mux_o_3572),
  .I0(ram16sdp_inst_263_dout[28]),
  .I1(ram16sdp_inst_271_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3573 (
  .O(mux_o_3573),
  .I0(ram16sdp_inst_279_dout[28]),
  .I1(ram16sdp_inst_287_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3574 (
  .O(mux_o_3574),
  .I0(ram16sdp_inst_295_dout[28]),
  .I1(ram16sdp_inst_303_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3575 (
  .O(mux_o_3575),
  .I0(ram16sdp_inst_311_dout[28]),
  .I1(ram16sdp_inst_319_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3576 (
  .O(mux_o_3576),
  .I0(ram16sdp_inst_327_dout[28]),
  .I1(ram16sdp_inst_335_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3577 (
  .O(mux_o_3577),
  .I0(ram16sdp_inst_343_dout[28]),
  .I1(ram16sdp_inst_351_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3578 (
  .O(mux_o_3578),
  .I0(ram16sdp_inst_359_dout[28]),
  .I1(ram16sdp_inst_367_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3579 (
  .O(mux_o_3579),
  .I0(ram16sdp_inst_375_dout[28]),
  .I1(ram16sdp_inst_383_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3580 (
  .O(mux_o_3580),
  .I0(ram16sdp_inst_391_dout[28]),
  .I1(ram16sdp_inst_399_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3581 (
  .O(mux_o_3581),
  .I0(ram16sdp_inst_407_dout[28]),
  .I1(ram16sdp_inst_415_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3582 (
  .O(mux_o_3582),
  .I0(ram16sdp_inst_423_dout[28]),
  .I1(ram16sdp_inst_431_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3583 (
  .O(mux_o_3583),
  .I0(ram16sdp_inst_439_dout[28]),
  .I1(ram16sdp_inst_447_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3584 (
  .O(mux_o_3584),
  .I0(ram16sdp_inst_455_dout[28]),
  .I1(ram16sdp_inst_463_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3585 (
  .O(mux_o_3585),
  .I0(ram16sdp_inst_471_dout[28]),
  .I1(ram16sdp_inst_479_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3586 (
  .O(mux_o_3586),
  .I0(ram16sdp_inst_487_dout[28]),
  .I1(ram16sdp_inst_495_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3587 (
  .O(mux_o_3587),
  .I0(ram16sdp_inst_503_dout[28]),
  .I1(ram16sdp_inst_511_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3588 (
  .O(mux_o_3588),
  .I0(ram16sdp_inst_519_dout[28]),
  .I1(ram16sdp_inst_527_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3589 (
  .O(mux_o_3589),
  .I0(ram16sdp_inst_535_dout[28]),
  .I1(ram16sdp_inst_543_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3590 (
  .O(mux_o_3590),
  .I0(ram16sdp_inst_551_dout[28]),
  .I1(ram16sdp_inst_559_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3591 (
  .O(mux_o_3591),
  .I0(ram16sdp_inst_567_dout[28]),
  .I1(ram16sdp_inst_575_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3592 (
  .O(mux_o_3592),
  .I0(ram16sdp_inst_583_dout[28]),
  .I1(ram16sdp_inst_591_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3593 (
  .O(mux_o_3593),
  .I0(ram16sdp_inst_599_dout[28]),
  .I1(ram16sdp_inst_607_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3594 (
  .O(mux_o_3594),
  .I0(ram16sdp_inst_615_dout[28]),
  .I1(ram16sdp_inst_623_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3595 (
  .O(mux_o_3595),
  .I0(ram16sdp_inst_631_dout[28]),
  .I1(ram16sdp_inst_639_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3596 (
  .O(mux_o_3596),
  .I0(ram16sdp_inst_647_dout[28]),
  .I1(ram16sdp_inst_655_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3597 (
  .O(mux_o_3597),
  .I0(ram16sdp_inst_663_dout[28]),
  .I1(ram16sdp_inst_671_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3598 (
  .O(mux_o_3598),
  .I0(ram16sdp_inst_679_dout[28]),
  .I1(ram16sdp_inst_687_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3599 (
  .O(mux_o_3599),
  .I0(ram16sdp_inst_695_dout[28]),
  .I1(ram16sdp_inst_703_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3600 (
  .O(mux_o_3600),
  .I0(ram16sdp_inst_711_dout[28]),
  .I1(ram16sdp_inst_719_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3601 (
  .O(mux_o_3601),
  .I0(ram16sdp_inst_727_dout[28]),
  .I1(ram16sdp_inst_735_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3602 (
  .O(mux_o_3602),
  .I0(ram16sdp_inst_743_dout[28]),
  .I1(ram16sdp_inst_751_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3603 (
  .O(mux_o_3603),
  .I0(ram16sdp_inst_759_dout[28]),
  .I1(ram16sdp_inst_767_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3604 (
  .O(mux_o_3604),
  .I0(ram16sdp_inst_775_dout[28]),
  .I1(ram16sdp_inst_783_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3605 (
  .O(mux_o_3605),
  .I0(ram16sdp_inst_791_dout[28]),
  .I1(ram16sdp_inst_799_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3606 (
  .O(mux_o_3606),
  .I0(ram16sdp_inst_807_dout[28]),
  .I1(ram16sdp_inst_815_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3607 (
  .O(mux_o_3607),
  .I0(ram16sdp_inst_823_dout[28]),
  .I1(ram16sdp_inst_831_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3608 (
  .O(mux_o_3608),
  .I0(ram16sdp_inst_839_dout[28]),
  .I1(ram16sdp_inst_847_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3609 (
  .O(mux_o_3609),
  .I0(ram16sdp_inst_855_dout[28]),
  .I1(ram16sdp_inst_863_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3610 (
  .O(mux_o_3610),
  .I0(ram16sdp_inst_871_dout[28]),
  .I1(ram16sdp_inst_879_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3611 (
  .O(mux_o_3611),
  .I0(ram16sdp_inst_887_dout[28]),
  .I1(ram16sdp_inst_895_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3612 (
  .O(mux_o_3612),
  .I0(ram16sdp_inst_903_dout[28]),
  .I1(ram16sdp_inst_911_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3613 (
  .O(mux_o_3613),
  .I0(ram16sdp_inst_919_dout[28]),
  .I1(ram16sdp_inst_927_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3614 (
  .O(mux_o_3614),
  .I0(ram16sdp_inst_935_dout[28]),
  .I1(ram16sdp_inst_943_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3615 (
  .O(mux_o_3615),
  .I0(ram16sdp_inst_951_dout[28]),
  .I1(ram16sdp_inst_959_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3616 (
  .O(mux_o_3616),
  .I0(ram16sdp_inst_967_dout[28]),
  .I1(ram16sdp_inst_975_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3617 (
  .O(mux_o_3617),
  .I0(ram16sdp_inst_983_dout[28]),
  .I1(ram16sdp_inst_991_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3618 (
  .O(mux_o_3618),
  .I0(ram16sdp_inst_999_dout[28]),
  .I1(ram16sdp_inst_1007_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3619 (
  .O(mux_o_3619),
  .I0(ram16sdp_inst_1015_dout[28]),
  .I1(ram16sdp_inst_1023_dout[28]),
  .S0(rad[4])
);
MUX2 mux_inst_3620 (
  .O(mux_o_3620),
  .I0(mux_o_3556),
  .I1(mux_o_3557),
  .S0(rad[5])
);
MUX2 mux_inst_3621 (
  .O(mux_o_3621),
  .I0(mux_o_3558),
  .I1(mux_o_3559),
  .S0(rad[5])
);
MUX2 mux_inst_3622 (
  .O(mux_o_3622),
  .I0(mux_o_3560),
  .I1(mux_o_3561),
  .S0(rad[5])
);
MUX2 mux_inst_3623 (
  .O(mux_o_3623),
  .I0(mux_o_3562),
  .I1(mux_o_3563),
  .S0(rad[5])
);
MUX2 mux_inst_3624 (
  .O(mux_o_3624),
  .I0(mux_o_3564),
  .I1(mux_o_3565),
  .S0(rad[5])
);
MUX2 mux_inst_3625 (
  .O(mux_o_3625),
  .I0(mux_o_3566),
  .I1(mux_o_3567),
  .S0(rad[5])
);
MUX2 mux_inst_3626 (
  .O(mux_o_3626),
  .I0(mux_o_3568),
  .I1(mux_o_3569),
  .S0(rad[5])
);
MUX2 mux_inst_3627 (
  .O(mux_o_3627),
  .I0(mux_o_3570),
  .I1(mux_o_3571),
  .S0(rad[5])
);
MUX2 mux_inst_3628 (
  .O(mux_o_3628),
  .I0(mux_o_3572),
  .I1(mux_o_3573),
  .S0(rad[5])
);
MUX2 mux_inst_3629 (
  .O(mux_o_3629),
  .I0(mux_o_3574),
  .I1(mux_o_3575),
  .S0(rad[5])
);
MUX2 mux_inst_3630 (
  .O(mux_o_3630),
  .I0(mux_o_3576),
  .I1(mux_o_3577),
  .S0(rad[5])
);
MUX2 mux_inst_3631 (
  .O(mux_o_3631),
  .I0(mux_o_3578),
  .I1(mux_o_3579),
  .S0(rad[5])
);
MUX2 mux_inst_3632 (
  .O(mux_o_3632),
  .I0(mux_o_3580),
  .I1(mux_o_3581),
  .S0(rad[5])
);
MUX2 mux_inst_3633 (
  .O(mux_o_3633),
  .I0(mux_o_3582),
  .I1(mux_o_3583),
  .S0(rad[5])
);
MUX2 mux_inst_3634 (
  .O(mux_o_3634),
  .I0(mux_o_3584),
  .I1(mux_o_3585),
  .S0(rad[5])
);
MUX2 mux_inst_3635 (
  .O(mux_o_3635),
  .I0(mux_o_3586),
  .I1(mux_o_3587),
  .S0(rad[5])
);
MUX2 mux_inst_3636 (
  .O(mux_o_3636),
  .I0(mux_o_3588),
  .I1(mux_o_3589),
  .S0(rad[5])
);
MUX2 mux_inst_3637 (
  .O(mux_o_3637),
  .I0(mux_o_3590),
  .I1(mux_o_3591),
  .S0(rad[5])
);
MUX2 mux_inst_3638 (
  .O(mux_o_3638),
  .I0(mux_o_3592),
  .I1(mux_o_3593),
  .S0(rad[5])
);
MUX2 mux_inst_3639 (
  .O(mux_o_3639),
  .I0(mux_o_3594),
  .I1(mux_o_3595),
  .S0(rad[5])
);
MUX2 mux_inst_3640 (
  .O(mux_o_3640),
  .I0(mux_o_3596),
  .I1(mux_o_3597),
  .S0(rad[5])
);
MUX2 mux_inst_3641 (
  .O(mux_o_3641),
  .I0(mux_o_3598),
  .I1(mux_o_3599),
  .S0(rad[5])
);
MUX2 mux_inst_3642 (
  .O(mux_o_3642),
  .I0(mux_o_3600),
  .I1(mux_o_3601),
  .S0(rad[5])
);
MUX2 mux_inst_3643 (
  .O(mux_o_3643),
  .I0(mux_o_3602),
  .I1(mux_o_3603),
  .S0(rad[5])
);
MUX2 mux_inst_3644 (
  .O(mux_o_3644),
  .I0(mux_o_3604),
  .I1(mux_o_3605),
  .S0(rad[5])
);
MUX2 mux_inst_3645 (
  .O(mux_o_3645),
  .I0(mux_o_3606),
  .I1(mux_o_3607),
  .S0(rad[5])
);
MUX2 mux_inst_3646 (
  .O(mux_o_3646),
  .I0(mux_o_3608),
  .I1(mux_o_3609),
  .S0(rad[5])
);
MUX2 mux_inst_3647 (
  .O(mux_o_3647),
  .I0(mux_o_3610),
  .I1(mux_o_3611),
  .S0(rad[5])
);
MUX2 mux_inst_3648 (
  .O(mux_o_3648),
  .I0(mux_o_3612),
  .I1(mux_o_3613),
  .S0(rad[5])
);
MUX2 mux_inst_3649 (
  .O(mux_o_3649),
  .I0(mux_o_3614),
  .I1(mux_o_3615),
  .S0(rad[5])
);
MUX2 mux_inst_3650 (
  .O(mux_o_3650),
  .I0(mux_o_3616),
  .I1(mux_o_3617),
  .S0(rad[5])
);
MUX2 mux_inst_3651 (
  .O(mux_o_3651),
  .I0(mux_o_3618),
  .I1(mux_o_3619),
  .S0(rad[5])
);
MUX2 mux_inst_3652 (
  .O(mux_o_3652),
  .I0(mux_o_3620),
  .I1(mux_o_3621),
  .S0(rad[6])
);
MUX2 mux_inst_3653 (
  .O(mux_o_3653),
  .I0(mux_o_3622),
  .I1(mux_o_3623),
  .S0(rad[6])
);
MUX2 mux_inst_3654 (
  .O(mux_o_3654),
  .I0(mux_o_3624),
  .I1(mux_o_3625),
  .S0(rad[6])
);
MUX2 mux_inst_3655 (
  .O(mux_o_3655),
  .I0(mux_o_3626),
  .I1(mux_o_3627),
  .S0(rad[6])
);
MUX2 mux_inst_3656 (
  .O(mux_o_3656),
  .I0(mux_o_3628),
  .I1(mux_o_3629),
  .S0(rad[6])
);
MUX2 mux_inst_3657 (
  .O(mux_o_3657),
  .I0(mux_o_3630),
  .I1(mux_o_3631),
  .S0(rad[6])
);
MUX2 mux_inst_3658 (
  .O(mux_o_3658),
  .I0(mux_o_3632),
  .I1(mux_o_3633),
  .S0(rad[6])
);
MUX2 mux_inst_3659 (
  .O(mux_o_3659),
  .I0(mux_o_3634),
  .I1(mux_o_3635),
  .S0(rad[6])
);
MUX2 mux_inst_3660 (
  .O(mux_o_3660),
  .I0(mux_o_3636),
  .I1(mux_o_3637),
  .S0(rad[6])
);
MUX2 mux_inst_3661 (
  .O(mux_o_3661),
  .I0(mux_o_3638),
  .I1(mux_o_3639),
  .S0(rad[6])
);
MUX2 mux_inst_3662 (
  .O(mux_o_3662),
  .I0(mux_o_3640),
  .I1(mux_o_3641),
  .S0(rad[6])
);
MUX2 mux_inst_3663 (
  .O(mux_o_3663),
  .I0(mux_o_3642),
  .I1(mux_o_3643),
  .S0(rad[6])
);
MUX2 mux_inst_3664 (
  .O(mux_o_3664),
  .I0(mux_o_3644),
  .I1(mux_o_3645),
  .S0(rad[6])
);
MUX2 mux_inst_3665 (
  .O(mux_o_3665),
  .I0(mux_o_3646),
  .I1(mux_o_3647),
  .S0(rad[6])
);
MUX2 mux_inst_3666 (
  .O(mux_o_3666),
  .I0(mux_o_3648),
  .I1(mux_o_3649),
  .S0(rad[6])
);
MUX2 mux_inst_3667 (
  .O(mux_o_3667),
  .I0(mux_o_3650),
  .I1(mux_o_3651),
  .S0(rad[6])
);
MUX2 mux_inst_3668 (
  .O(mux_o_3668),
  .I0(mux_o_3652),
  .I1(mux_o_3653),
  .S0(rad[7])
);
MUX2 mux_inst_3669 (
  .O(mux_o_3669),
  .I0(mux_o_3654),
  .I1(mux_o_3655),
  .S0(rad[7])
);
MUX2 mux_inst_3670 (
  .O(mux_o_3670),
  .I0(mux_o_3656),
  .I1(mux_o_3657),
  .S0(rad[7])
);
MUX2 mux_inst_3671 (
  .O(mux_o_3671),
  .I0(mux_o_3658),
  .I1(mux_o_3659),
  .S0(rad[7])
);
MUX2 mux_inst_3672 (
  .O(mux_o_3672),
  .I0(mux_o_3660),
  .I1(mux_o_3661),
  .S0(rad[7])
);
MUX2 mux_inst_3673 (
  .O(mux_o_3673),
  .I0(mux_o_3662),
  .I1(mux_o_3663),
  .S0(rad[7])
);
MUX2 mux_inst_3674 (
  .O(mux_o_3674),
  .I0(mux_o_3664),
  .I1(mux_o_3665),
  .S0(rad[7])
);
MUX2 mux_inst_3675 (
  .O(mux_o_3675),
  .I0(mux_o_3666),
  .I1(mux_o_3667),
  .S0(rad[7])
);
MUX2 mux_inst_3676 (
  .O(mux_o_3676),
  .I0(mux_o_3668),
  .I1(mux_o_3669),
  .S0(rad[8])
);
MUX2 mux_inst_3677 (
  .O(mux_o_3677),
  .I0(mux_o_3670),
  .I1(mux_o_3671),
  .S0(rad[8])
);
MUX2 mux_inst_3678 (
  .O(mux_o_3678),
  .I0(mux_o_3672),
  .I1(mux_o_3673),
  .S0(rad[8])
);
MUX2 mux_inst_3679 (
  .O(mux_o_3679),
  .I0(mux_o_3674),
  .I1(mux_o_3675),
  .S0(rad[8])
);
MUX2 mux_inst_3680 (
  .O(mux_o_3680),
  .I0(mux_o_3676),
  .I1(mux_o_3677),
  .S0(rad[9])
);
MUX2 mux_inst_3681 (
  .O(mux_o_3681),
  .I0(mux_o_3678),
  .I1(mux_o_3679),
  .S0(rad[9])
);
MUX2 mux_inst_3682 (
  .O(dout[28]),
  .I0(mux_o_3680),
  .I1(mux_o_3681),
  .S0(rad[10])
);
MUX2 mux_inst_3683 (
  .O(mux_o_3683),
  .I0(ram16sdp_inst_7_dout[29]),
  .I1(ram16sdp_inst_15_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3684 (
  .O(mux_o_3684),
  .I0(ram16sdp_inst_23_dout[29]),
  .I1(ram16sdp_inst_31_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3685 (
  .O(mux_o_3685),
  .I0(ram16sdp_inst_39_dout[29]),
  .I1(ram16sdp_inst_47_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3686 (
  .O(mux_o_3686),
  .I0(ram16sdp_inst_55_dout[29]),
  .I1(ram16sdp_inst_63_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3687 (
  .O(mux_o_3687),
  .I0(ram16sdp_inst_71_dout[29]),
  .I1(ram16sdp_inst_79_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3688 (
  .O(mux_o_3688),
  .I0(ram16sdp_inst_87_dout[29]),
  .I1(ram16sdp_inst_95_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3689 (
  .O(mux_o_3689),
  .I0(ram16sdp_inst_103_dout[29]),
  .I1(ram16sdp_inst_111_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3690 (
  .O(mux_o_3690),
  .I0(ram16sdp_inst_119_dout[29]),
  .I1(ram16sdp_inst_127_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3691 (
  .O(mux_o_3691),
  .I0(ram16sdp_inst_135_dout[29]),
  .I1(ram16sdp_inst_143_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3692 (
  .O(mux_o_3692),
  .I0(ram16sdp_inst_151_dout[29]),
  .I1(ram16sdp_inst_159_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3693 (
  .O(mux_o_3693),
  .I0(ram16sdp_inst_167_dout[29]),
  .I1(ram16sdp_inst_175_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3694 (
  .O(mux_o_3694),
  .I0(ram16sdp_inst_183_dout[29]),
  .I1(ram16sdp_inst_191_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3695 (
  .O(mux_o_3695),
  .I0(ram16sdp_inst_199_dout[29]),
  .I1(ram16sdp_inst_207_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3696 (
  .O(mux_o_3696),
  .I0(ram16sdp_inst_215_dout[29]),
  .I1(ram16sdp_inst_223_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3697 (
  .O(mux_o_3697),
  .I0(ram16sdp_inst_231_dout[29]),
  .I1(ram16sdp_inst_239_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3698 (
  .O(mux_o_3698),
  .I0(ram16sdp_inst_247_dout[29]),
  .I1(ram16sdp_inst_255_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3699 (
  .O(mux_o_3699),
  .I0(ram16sdp_inst_263_dout[29]),
  .I1(ram16sdp_inst_271_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3700 (
  .O(mux_o_3700),
  .I0(ram16sdp_inst_279_dout[29]),
  .I1(ram16sdp_inst_287_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3701 (
  .O(mux_o_3701),
  .I0(ram16sdp_inst_295_dout[29]),
  .I1(ram16sdp_inst_303_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3702 (
  .O(mux_o_3702),
  .I0(ram16sdp_inst_311_dout[29]),
  .I1(ram16sdp_inst_319_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3703 (
  .O(mux_o_3703),
  .I0(ram16sdp_inst_327_dout[29]),
  .I1(ram16sdp_inst_335_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3704 (
  .O(mux_o_3704),
  .I0(ram16sdp_inst_343_dout[29]),
  .I1(ram16sdp_inst_351_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3705 (
  .O(mux_o_3705),
  .I0(ram16sdp_inst_359_dout[29]),
  .I1(ram16sdp_inst_367_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3706 (
  .O(mux_o_3706),
  .I0(ram16sdp_inst_375_dout[29]),
  .I1(ram16sdp_inst_383_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3707 (
  .O(mux_o_3707),
  .I0(ram16sdp_inst_391_dout[29]),
  .I1(ram16sdp_inst_399_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3708 (
  .O(mux_o_3708),
  .I0(ram16sdp_inst_407_dout[29]),
  .I1(ram16sdp_inst_415_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3709 (
  .O(mux_o_3709),
  .I0(ram16sdp_inst_423_dout[29]),
  .I1(ram16sdp_inst_431_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3710 (
  .O(mux_o_3710),
  .I0(ram16sdp_inst_439_dout[29]),
  .I1(ram16sdp_inst_447_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3711 (
  .O(mux_o_3711),
  .I0(ram16sdp_inst_455_dout[29]),
  .I1(ram16sdp_inst_463_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3712 (
  .O(mux_o_3712),
  .I0(ram16sdp_inst_471_dout[29]),
  .I1(ram16sdp_inst_479_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3713 (
  .O(mux_o_3713),
  .I0(ram16sdp_inst_487_dout[29]),
  .I1(ram16sdp_inst_495_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3714 (
  .O(mux_o_3714),
  .I0(ram16sdp_inst_503_dout[29]),
  .I1(ram16sdp_inst_511_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3715 (
  .O(mux_o_3715),
  .I0(ram16sdp_inst_519_dout[29]),
  .I1(ram16sdp_inst_527_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3716 (
  .O(mux_o_3716),
  .I0(ram16sdp_inst_535_dout[29]),
  .I1(ram16sdp_inst_543_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3717 (
  .O(mux_o_3717),
  .I0(ram16sdp_inst_551_dout[29]),
  .I1(ram16sdp_inst_559_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3718 (
  .O(mux_o_3718),
  .I0(ram16sdp_inst_567_dout[29]),
  .I1(ram16sdp_inst_575_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3719 (
  .O(mux_o_3719),
  .I0(ram16sdp_inst_583_dout[29]),
  .I1(ram16sdp_inst_591_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3720 (
  .O(mux_o_3720),
  .I0(ram16sdp_inst_599_dout[29]),
  .I1(ram16sdp_inst_607_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3721 (
  .O(mux_o_3721),
  .I0(ram16sdp_inst_615_dout[29]),
  .I1(ram16sdp_inst_623_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3722 (
  .O(mux_o_3722),
  .I0(ram16sdp_inst_631_dout[29]),
  .I1(ram16sdp_inst_639_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3723 (
  .O(mux_o_3723),
  .I0(ram16sdp_inst_647_dout[29]),
  .I1(ram16sdp_inst_655_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3724 (
  .O(mux_o_3724),
  .I0(ram16sdp_inst_663_dout[29]),
  .I1(ram16sdp_inst_671_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3725 (
  .O(mux_o_3725),
  .I0(ram16sdp_inst_679_dout[29]),
  .I1(ram16sdp_inst_687_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3726 (
  .O(mux_o_3726),
  .I0(ram16sdp_inst_695_dout[29]),
  .I1(ram16sdp_inst_703_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3727 (
  .O(mux_o_3727),
  .I0(ram16sdp_inst_711_dout[29]),
  .I1(ram16sdp_inst_719_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3728 (
  .O(mux_o_3728),
  .I0(ram16sdp_inst_727_dout[29]),
  .I1(ram16sdp_inst_735_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3729 (
  .O(mux_o_3729),
  .I0(ram16sdp_inst_743_dout[29]),
  .I1(ram16sdp_inst_751_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3730 (
  .O(mux_o_3730),
  .I0(ram16sdp_inst_759_dout[29]),
  .I1(ram16sdp_inst_767_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3731 (
  .O(mux_o_3731),
  .I0(ram16sdp_inst_775_dout[29]),
  .I1(ram16sdp_inst_783_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3732 (
  .O(mux_o_3732),
  .I0(ram16sdp_inst_791_dout[29]),
  .I1(ram16sdp_inst_799_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3733 (
  .O(mux_o_3733),
  .I0(ram16sdp_inst_807_dout[29]),
  .I1(ram16sdp_inst_815_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3734 (
  .O(mux_o_3734),
  .I0(ram16sdp_inst_823_dout[29]),
  .I1(ram16sdp_inst_831_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3735 (
  .O(mux_o_3735),
  .I0(ram16sdp_inst_839_dout[29]),
  .I1(ram16sdp_inst_847_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3736 (
  .O(mux_o_3736),
  .I0(ram16sdp_inst_855_dout[29]),
  .I1(ram16sdp_inst_863_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3737 (
  .O(mux_o_3737),
  .I0(ram16sdp_inst_871_dout[29]),
  .I1(ram16sdp_inst_879_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3738 (
  .O(mux_o_3738),
  .I0(ram16sdp_inst_887_dout[29]),
  .I1(ram16sdp_inst_895_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3739 (
  .O(mux_o_3739),
  .I0(ram16sdp_inst_903_dout[29]),
  .I1(ram16sdp_inst_911_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3740 (
  .O(mux_o_3740),
  .I0(ram16sdp_inst_919_dout[29]),
  .I1(ram16sdp_inst_927_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3741 (
  .O(mux_o_3741),
  .I0(ram16sdp_inst_935_dout[29]),
  .I1(ram16sdp_inst_943_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3742 (
  .O(mux_o_3742),
  .I0(ram16sdp_inst_951_dout[29]),
  .I1(ram16sdp_inst_959_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3743 (
  .O(mux_o_3743),
  .I0(ram16sdp_inst_967_dout[29]),
  .I1(ram16sdp_inst_975_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3744 (
  .O(mux_o_3744),
  .I0(ram16sdp_inst_983_dout[29]),
  .I1(ram16sdp_inst_991_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3745 (
  .O(mux_o_3745),
  .I0(ram16sdp_inst_999_dout[29]),
  .I1(ram16sdp_inst_1007_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3746 (
  .O(mux_o_3746),
  .I0(ram16sdp_inst_1015_dout[29]),
  .I1(ram16sdp_inst_1023_dout[29]),
  .S0(rad[4])
);
MUX2 mux_inst_3747 (
  .O(mux_o_3747),
  .I0(mux_o_3683),
  .I1(mux_o_3684),
  .S0(rad[5])
);
MUX2 mux_inst_3748 (
  .O(mux_o_3748),
  .I0(mux_o_3685),
  .I1(mux_o_3686),
  .S0(rad[5])
);
MUX2 mux_inst_3749 (
  .O(mux_o_3749),
  .I0(mux_o_3687),
  .I1(mux_o_3688),
  .S0(rad[5])
);
MUX2 mux_inst_3750 (
  .O(mux_o_3750),
  .I0(mux_o_3689),
  .I1(mux_o_3690),
  .S0(rad[5])
);
MUX2 mux_inst_3751 (
  .O(mux_o_3751),
  .I0(mux_o_3691),
  .I1(mux_o_3692),
  .S0(rad[5])
);
MUX2 mux_inst_3752 (
  .O(mux_o_3752),
  .I0(mux_o_3693),
  .I1(mux_o_3694),
  .S0(rad[5])
);
MUX2 mux_inst_3753 (
  .O(mux_o_3753),
  .I0(mux_o_3695),
  .I1(mux_o_3696),
  .S0(rad[5])
);
MUX2 mux_inst_3754 (
  .O(mux_o_3754),
  .I0(mux_o_3697),
  .I1(mux_o_3698),
  .S0(rad[5])
);
MUX2 mux_inst_3755 (
  .O(mux_o_3755),
  .I0(mux_o_3699),
  .I1(mux_o_3700),
  .S0(rad[5])
);
MUX2 mux_inst_3756 (
  .O(mux_o_3756),
  .I0(mux_o_3701),
  .I1(mux_o_3702),
  .S0(rad[5])
);
MUX2 mux_inst_3757 (
  .O(mux_o_3757),
  .I0(mux_o_3703),
  .I1(mux_o_3704),
  .S0(rad[5])
);
MUX2 mux_inst_3758 (
  .O(mux_o_3758),
  .I0(mux_o_3705),
  .I1(mux_o_3706),
  .S0(rad[5])
);
MUX2 mux_inst_3759 (
  .O(mux_o_3759),
  .I0(mux_o_3707),
  .I1(mux_o_3708),
  .S0(rad[5])
);
MUX2 mux_inst_3760 (
  .O(mux_o_3760),
  .I0(mux_o_3709),
  .I1(mux_o_3710),
  .S0(rad[5])
);
MUX2 mux_inst_3761 (
  .O(mux_o_3761),
  .I0(mux_o_3711),
  .I1(mux_o_3712),
  .S0(rad[5])
);
MUX2 mux_inst_3762 (
  .O(mux_o_3762),
  .I0(mux_o_3713),
  .I1(mux_o_3714),
  .S0(rad[5])
);
MUX2 mux_inst_3763 (
  .O(mux_o_3763),
  .I0(mux_o_3715),
  .I1(mux_o_3716),
  .S0(rad[5])
);
MUX2 mux_inst_3764 (
  .O(mux_o_3764),
  .I0(mux_o_3717),
  .I1(mux_o_3718),
  .S0(rad[5])
);
MUX2 mux_inst_3765 (
  .O(mux_o_3765),
  .I0(mux_o_3719),
  .I1(mux_o_3720),
  .S0(rad[5])
);
MUX2 mux_inst_3766 (
  .O(mux_o_3766),
  .I0(mux_o_3721),
  .I1(mux_o_3722),
  .S0(rad[5])
);
MUX2 mux_inst_3767 (
  .O(mux_o_3767),
  .I0(mux_o_3723),
  .I1(mux_o_3724),
  .S0(rad[5])
);
MUX2 mux_inst_3768 (
  .O(mux_o_3768),
  .I0(mux_o_3725),
  .I1(mux_o_3726),
  .S0(rad[5])
);
MUX2 mux_inst_3769 (
  .O(mux_o_3769),
  .I0(mux_o_3727),
  .I1(mux_o_3728),
  .S0(rad[5])
);
MUX2 mux_inst_3770 (
  .O(mux_o_3770),
  .I0(mux_o_3729),
  .I1(mux_o_3730),
  .S0(rad[5])
);
MUX2 mux_inst_3771 (
  .O(mux_o_3771),
  .I0(mux_o_3731),
  .I1(mux_o_3732),
  .S0(rad[5])
);
MUX2 mux_inst_3772 (
  .O(mux_o_3772),
  .I0(mux_o_3733),
  .I1(mux_o_3734),
  .S0(rad[5])
);
MUX2 mux_inst_3773 (
  .O(mux_o_3773),
  .I0(mux_o_3735),
  .I1(mux_o_3736),
  .S0(rad[5])
);
MUX2 mux_inst_3774 (
  .O(mux_o_3774),
  .I0(mux_o_3737),
  .I1(mux_o_3738),
  .S0(rad[5])
);
MUX2 mux_inst_3775 (
  .O(mux_o_3775),
  .I0(mux_o_3739),
  .I1(mux_o_3740),
  .S0(rad[5])
);
MUX2 mux_inst_3776 (
  .O(mux_o_3776),
  .I0(mux_o_3741),
  .I1(mux_o_3742),
  .S0(rad[5])
);
MUX2 mux_inst_3777 (
  .O(mux_o_3777),
  .I0(mux_o_3743),
  .I1(mux_o_3744),
  .S0(rad[5])
);
MUX2 mux_inst_3778 (
  .O(mux_o_3778),
  .I0(mux_o_3745),
  .I1(mux_o_3746),
  .S0(rad[5])
);
MUX2 mux_inst_3779 (
  .O(mux_o_3779),
  .I0(mux_o_3747),
  .I1(mux_o_3748),
  .S0(rad[6])
);
MUX2 mux_inst_3780 (
  .O(mux_o_3780),
  .I0(mux_o_3749),
  .I1(mux_o_3750),
  .S0(rad[6])
);
MUX2 mux_inst_3781 (
  .O(mux_o_3781),
  .I0(mux_o_3751),
  .I1(mux_o_3752),
  .S0(rad[6])
);
MUX2 mux_inst_3782 (
  .O(mux_o_3782),
  .I0(mux_o_3753),
  .I1(mux_o_3754),
  .S0(rad[6])
);
MUX2 mux_inst_3783 (
  .O(mux_o_3783),
  .I0(mux_o_3755),
  .I1(mux_o_3756),
  .S0(rad[6])
);
MUX2 mux_inst_3784 (
  .O(mux_o_3784),
  .I0(mux_o_3757),
  .I1(mux_o_3758),
  .S0(rad[6])
);
MUX2 mux_inst_3785 (
  .O(mux_o_3785),
  .I0(mux_o_3759),
  .I1(mux_o_3760),
  .S0(rad[6])
);
MUX2 mux_inst_3786 (
  .O(mux_o_3786),
  .I0(mux_o_3761),
  .I1(mux_o_3762),
  .S0(rad[6])
);
MUX2 mux_inst_3787 (
  .O(mux_o_3787),
  .I0(mux_o_3763),
  .I1(mux_o_3764),
  .S0(rad[6])
);
MUX2 mux_inst_3788 (
  .O(mux_o_3788),
  .I0(mux_o_3765),
  .I1(mux_o_3766),
  .S0(rad[6])
);
MUX2 mux_inst_3789 (
  .O(mux_o_3789),
  .I0(mux_o_3767),
  .I1(mux_o_3768),
  .S0(rad[6])
);
MUX2 mux_inst_3790 (
  .O(mux_o_3790),
  .I0(mux_o_3769),
  .I1(mux_o_3770),
  .S0(rad[6])
);
MUX2 mux_inst_3791 (
  .O(mux_o_3791),
  .I0(mux_o_3771),
  .I1(mux_o_3772),
  .S0(rad[6])
);
MUX2 mux_inst_3792 (
  .O(mux_o_3792),
  .I0(mux_o_3773),
  .I1(mux_o_3774),
  .S0(rad[6])
);
MUX2 mux_inst_3793 (
  .O(mux_o_3793),
  .I0(mux_o_3775),
  .I1(mux_o_3776),
  .S0(rad[6])
);
MUX2 mux_inst_3794 (
  .O(mux_o_3794),
  .I0(mux_o_3777),
  .I1(mux_o_3778),
  .S0(rad[6])
);
MUX2 mux_inst_3795 (
  .O(mux_o_3795),
  .I0(mux_o_3779),
  .I1(mux_o_3780),
  .S0(rad[7])
);
MUX2 mux_inst_3796 (
  .O(mux_o_3796),
  .I0(mux_o_3781),
  .I1(mux_o_3782),
  .S0(rad[7])
);
MUX2 mux_inst_3797 (
  .O(mux_o_3797),
  .I0(mux_o_3783),
  .I1(mux_o_3784),
  .S0(rad[7])
);
MUX2 mux_inst_3798 (
  .O(mux_o_3798),
  .I0(mux_o_3785),
  .I1(mux_o_3786),
  .S0(rad[7])
);
MUX2 mux_inst_3799 (
  .O(mux_o_3799),
  .I0(mux_o_3787),
  .I1(mux_o_3788),
  .S0(rad[7])
);
MUX2 mux_inst_3800 (
  .O(mux_o_3800),
  .I0(mux_o_3789),
  .I1(mux_o_3790),
  .S0(rad[7])
);
MUX2 mux_inst_3801 (
  .O(mux_o_3801),
  .I0(mux_o_3791),
  .I1(mux_o_3792),
  .S0(rad[7])
);
MUX2 mux_inst_3802 (
  .O(mux_o_3802),
  .I0(mux_o_3793),
  .I1(mux_o_3794),
  .S0(rad[7])
);
MUX2 mux_inst_3803 (
  .O(mux_o_3803),
  .I0(mux_o_3795),
  .I1(mux_o_3796),
  .S0(rad[8])
);
MUX2 mux_inst_3804 (
  .O(mux_o_3804),
  .I0(mux_o_3797),
  .I1(mux_o_3798),
  .S0(rad[8])
);
MUX2 mux_inst_3805 (
  .O(mux_o_3805),
  .I0(mux_o_3799),
  .I1(mux_o_3800),
  .S0(rad[8])
);
MUX2 mux_inst_3806 (
  .O(mux_o_3806),
  .I0(mux_o_3801),
  .I1(mux_o_3802),
  .S0(rad[8])
);
MUX2 mux_inst_3807 (
  .O(mux_o_3807),
  .I0(mux_o_3803),
  .I1(mux_o_3804),
  .S0(rad[9])
);
MUX2 mux_inst_3808 (
  .O(mux_o_3808),
  .I0(mux_o_3805),
  .I1(mux_o_3806),
  .S0(rad[9])
);
MUX2 mux_inst_3809 (
  .O(dout[29]),
  .I0(mux_o_3807),
  .I1(mux_o_3808),
  .S0(rad[10])
);
MUX2 mux_inst_3810 (
  .O(mux_o_3810),
  .I0(ram16sdp_inst_7_dout[30]),
  .I1(ram16sdp_inst_15_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3811 (
  .O(mux_o_3811),
  .I0(ram16sdp_inst_23_dout[30]),
  .I1(ram16sdp_inst_31_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3812 (
  .O(mux_o_3812),
  .I0(ram16sdp_inst_39_dout[30]),
  .I1(ram16sdp_inst_47_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3813 (
  .O(mux_o_3813),
  .I0(ram16sdp_inst_55_dout[30]),
  .I1(ram16sdp_inst_63_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3814 (
  .O(mux_o_3814),
  .I0(ram16sdp_inst_71_dout[30]),
  .I1(ram16sdp_inst_79_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3815 (
  .O(mux_o_3815),
  .I0(ram16sdp_inst_87_dout[30]),
  .I1(ram16sdp_inst_95_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3816 (
  .O(mux_o_3816),
  .I0(ram16sdp_inst_103_dout[30]),
  .I1(ram16sdp_inst_111_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3817 (
  .O(mux_o_3817),
  .I0(ram16sdp_inst_119_dout[30]),
  .I1(ram16sdp_inst_127_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3818 (
  .O(mux_o_3818),
  .I0(ram16sdp_inst_135_dout[30]),
  .I1(ram16sdp_inst_143_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3819 (
  .O(mux_o_3819),
  .I0(ram16sdp_inst_151_dout[30]),
  .I1(ram16sdp_inst_159_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3820 (
  .O(mux_o_3820),
  .I0(ram16sdp_inst_167_dout[30]),
  .I1(ram16sdp_inst_175_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3821 (
  .O(mux_o_3821),
  .I0(ram16sdp_inst_183_dout[30]),
  .I1(ram16sdp_inst_191_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3822 (
  .O(mux_o_3822),
  .I0(ram16sdp_inst_199_dout[30]),
  .I1(ram16sdp_inst_207_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3823 (
  .O(mux_o_3823),
  .I0(ram16sdp_inst_215_dout[30]),
  .I1(ram16sdp_inst_223_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3824 (
  .O(mux_o_3824),
  .I0(ram16sdp_inst_231_dout[30]),
  .I1(ram16sdp_inst_239_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3825 (
  .O(mux_o_3825),
  .I0(ram16sdp_inst_247_dout[30]),
  .I1(ram16sdp_inst_255_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3826 (
  .O(mux_o_3826),
  .I0(ram16sdp_inst_263_dout[30]),
  .I1(ram16sdp_inst_271_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3827 (
  .O(mux_o_3827),
  .I0(ram16sdp_inst_279_dout[30]),
  .I1(ram16sdp_inst_287_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3828 (
  .O(mux_o_3828),
  .I0(ram16sdp_inst_295_dout[30]),
  .I1(ram16sdp_inst_303_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3829 (
  .O(mux_o_3829),
  .I0(ram16sdp_inst_311_dout[30]),
  .I1(ram16sdp_inst_319_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3830 (
  .O(mux_o_3830),
  .I0(ram16sdp_inst_327_dout[30]),
  .I1(ram16sdp_inst_335_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3831 (
  .O(mux_o_3831),
  .I0(ram16sdp_inst_343_dout[30]),
  .I1(ram16sdp_inst_351_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3832 (
  .O(mux_o_3832),
  .I0(ram16sdp_inst_359_dout[30]),
  .I1(ram16sdp_inst_367_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3833 (
  .O(mux_o_3833),
  .I0(ram16sdp_inst_375_dout[30]),
  .I1(ram16sdp_inst_383_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3834 (
  .O(mux_o_3834),
  .I0(ram16sdp_inst_391_dout[30]),
  .I1(ram16sdp_inst_399_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3835 (
  .O(mux_o_3835),
  .I0(ram16sdp_inst_407_dout[30]),
  .I1(ram16sdp_inst_415_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3836 (
  .O(mux_o_3836),
  .I0(ram16sdp_inst_423_dout[30]),
  .I1(ram16sdp_inst_431_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3837 (
  .O(mux_o_3837),
  .I0(ram16sdp_inst_439_dout[30]),
  .I1(ram16sdp_inst_447_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3838 (
  .O(mux_o_3838),
  .I0(ram16sdp_inst_455_dout[30]),
  .I1(ram16sdp_inst_463_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3839 (
  .O(mux_o_3839),
  .I0(ram16sdp_inst_471_dout[30]),
  .I1(ram16sdp_inst_479_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3840 (
  .O(mux_o_3840),
  .I0(ram16sdp_inst_487_dout[30]),
  .I1(ram16sdp_inst_495_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3841 (
  .O(mux_o_3841),
  .I0(ram16sdp_inst_503_dout[30]),
  .I1(ram16sdp_inst_511_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3842 (
  .O(mux_o_3842),
  .I0(ram16sdp_inst_519_dout[30]),
  .I1(ram16sdp_inst_527_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3843 (
  .O(mux_o_3843),
  .I0(ram16sdp_inst_535_dout[30]),
  .I1(ram16sdp_inst_543_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3844 (
  .O(mux_o_3844),
  .I0(ram16sdp_inst_551_dout[30]),
  .I1(ram16sdp_inst_559_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3845 (
  .O(mux_o_3845),
  .I0(ram16sdp_inst_567_dout[30]),
  .I1(ram16sdp_inst_575_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3846 (
  .O(mux_o_3846),
  .I0(ram16sdp_inst_583_dout[30]),
  .I1(ram16sdp_inst_591_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3847 (
  .O(mux_o_3847),
  .I0(ram16sdp_inst_599_dout[30]),
  .I1(ram16sdp_inst_607_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3848 (
  .O(mux_o_3848),
  .I0(ram16sdp_inst_615_dout[30]),
  .I1(ram16sdp_inst_623_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3849 (
  .O(mux_o_3849),
  .I0(ram16sdp_inst_631_dout[30]),
  .I1(ram16sdp_inst_639_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3850 (
  .O(mux_o_3850),
  .I0(ram16sdp_inst_647_dout[30]),
  .I1(ram16sdp_inst_655_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3851 (
  .O(mux_o_3851),
  .I0(ram16sdp_inst_663_dout[30]),
  .I1(ram16sdp_inst_671_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3852 (
  .O(mux_o_3852),
  .I0(ram16sdp_inst_679_dout[30]),
  .I1(ram16sdp_inst_687_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3853 (
  .O(mux_o_3853),
  .I0(ram16sdp_inst_695_dout[30]),
  .I1(ram16sdp_inst_703_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3854 (
  .O(mux_o_3854),
  .I0(ram16sdp_inst_711_dout[30]),
  .I1(ram16sdp_inst_719_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3855 (
  .O(mux_o_3855),
  .I0(ram16sdp_inst_727_dout[30]),
  .I1(ram16sdp_inst_735_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3856 (
  .O(mux_o_3856),
  .I0(ram16sdp_inst_743_dout[30]),
  .I1(ram16sdp_inst_751_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3857 (
  .O(mux_o_3857),
  .I0(ram16sdp_inst_759_dout[30]),
  .I1(ram16sdp_inst_767_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3858 (
  .O(mux_o_3858),
  .I0(ram16sdp_inst_775_dout[30]),
  .I1(ram16sdp_inst_783_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3859 (
  .O(mux_o_3859),
  .I0(ram16sdp_inst_791_dout[30]),
  .I1(ram16sdp_inst_799_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3860 (
  .O(mux_o_3860),
  .I0(ram16sdp_inst_807_dout[30]),
  .I1(ram16sdp_inst_815_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3861 (
  .O(mux_o_3861),
  .I0(ram16sdp_inst_823_dout[30]),
  .I1(ram16sdp_inst_831_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3862 (
  .O(mux_o_3862),
  .I0(ram16sdp_inst_839_dout[30]),
  .I1(ram16sdp_inst_847_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3863 (
  .O(mux_o_3863),
  .I0(ram16sdp_inst_855_dout[30]),
  .I1(ram16sdp_inst_863_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3864 (
  .O(mux_o_3864),
  .I0(ram16sdp_inst_871_dout[30]),
  .I1(ram16sdp_inst_879_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3865 (
  .O(mux_o_3865),
  .I0(ram16sdp_inst_887_dout[30]),
  .I1(ram16sdp_inst_895_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3866 (
  .O(mux_o_3866),
  .I0(ram16sdp_inst_903_dout[30]),
  .I1(ram16sdp_inst_911_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3867 (
  .O(mux_o_3867),
  .I0(ram16sdp_inst_919_dout[30]),
  .I1(ram16sdp_inst_927_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3868 (
  .O(mux_o_3868),
  .I0(ram16sdp_inst_935_dout[30]),
  .I1(ram16sdp_inst_943_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3869 (
  .O(mux_o_3869),
  .I0(ram16sdp_inst_951_dout[30]),
  .I1(ram16sdp_inst_959_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3870 (
  .O(mux_o_3870),
  .I0(ram16sdp_inst_967_dout[30]),
  .I1(ram16sdp_inst_975_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3871 (
  .O(mux_o_3871),
  .I0(ram16sdp_inst_983_dout[30]),
  .I1(ram16sdp_inst_991_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3872 (
  .O(mux_o_3872),
  .I0(ram16sdp_inst_999_dout[30]),
  .I1(ram16sdp_inst_1007_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3873 (
  .O(mux_o_3873),
  .I0(ram16sdp_inst_1015_dout[30]),
  .I1(ram16sdp_inst_1023_dout[30]),
  .S0(rad[4])
);
MUX2 mux_inst_3874 (
  .O(mux_o_3874),
  .I0(mux_o_3810),
  .I1(mux_o_3811),
  .S0(rad[5])
);
MUX2 mux_inst_3875 (
  .O(mux_o_3875),
  .I0(mux_o_3812),
  .I1(mux_o_3813),
  .S0(rad[5])
);
MUX2 mux_inst_3876 (
  .O(mux_o_3876),
  .I0(mux_o_3814),
  .I1(mux_o_3815),
  .S0(rad[5])
);
MUX2 mux_inst_3877 (
  .O(mux_o_3877),
  .I0(mux_o_3816),
  .I1(mux_o_3817),
  .S0(rad[5])
);
MUX2 mux_inst_3878 (
  .O(mux_o_3878),
  .I0(mux_o_3818),
  .I1(mux_o_3819),
  .S0(rad[5])
);
MUX2 mux_inst_3879 (
  .O(mux_o_3879),
  .I0(mux_o_3820),
  .I1(mux_o_3821),
  .S0(rad[5])
);
MUX2 mux_inst_3880 (
  .O(mux_o_3880),
  .I0(mux_o_3822),
  .I1(mux_o_3823),
  .S0(rad[5])
);
MUX2 mux_inst_3881 (
  .O(mux_o_3881),
  .I0(mux_o_3824),
  .I1(mux_o_3825),
  .S0(rad[5])
);
MUX2 mux_inst_3882 (
  .O(mux_o_3882),
  .I0(mux_o_3826),
  .I1(mux_o_3827),
  .S0(rad[5])
);
MUX2 mux_inst_3883 (
  .O(mux_o_3883),
  .I0(mux_o_3828),
  .I1(mux_o_3829),
  .S0(rad[5])
);
MUX2 mux_inst_3884 (
  .O(mux_o_3884),
  .I0(mux_o_3830),
  .I1(mux_o_3831),
  .S0(rad[5])
);
MUX2 mux_inst_3885 (
  .O(mux_o_3885),
  .I0(mux_o_3832),
  .I1(mux_o_3833),
  .S0(rad[5])
);
MUX2 mux_inst_3886 (
  .O(mux_o_3886),
  .I0(mux_o_3834),
  .I1(mux_o_3835),
  .S0(rad[5])
);
MUX2 mux_inst_3887 (
  .O(mux_o_3887),
  .I0(mux_o_3836),
  .I1(mux_o_3837),
  .S0(rad[5])
);
MUX2 mux_inst_3888 (
  .O(mux_o_3888),
  .I0(mux_o_3838),
  .I1(mux_o_3839),
  .S0(rad[5])
);
MUX2 mux_inst_3889 (
  .O(mux_o_3889),
  .I0(mux_o_3840),
  .I1(mux_o_3841),
  .S0(rad[5])
);
MUX2 mux_inst_3890 (
  .O(mux_o_3890),
  .I0(mux_o_3842),
  .I1(mux_o_3843),
  .S0(rad[5])
);
MUX2 mux_inst_3891 (
  .O(mux_o_3891),
  .I0(mux_o_3844),
  .I1(mux_o_3845),
  .S0(rad[5])
);
MUX2 mux_inst_3892 (
  .O(mux_o_3892),
  .I0(mux_o_3846),
  .I1(mux_o_3847),
  .S0(rad[5])
);
MUX2 mux_inst_3893 (
  .O(mux_o_3893),
  .I0(mux_o_3848),
  .I1(mux_o_3849),
  .S0(rad[5])
);
MUX2 mux_inst_3894 (
  .O(mux_o_3894),
  .I0(mux_o_3850),
  .I1(mux_o_3851),
  .S0(rad[5])
);
MUX2 mux_inst_3895 (
  .O(mux_o_3895),
  .I0(mux_o_3852),
  .I1(mux_o_3853),
  .S0(rad[5])
);
MUX2 mux_inst_3896 (
  .O(mux_o_3896),
  .I0(mux_o_3854),
  .I1(mux_o_3855),
  .S0(rad[5])
);
MUX2 mux_inst_3897 (
  .O(mux_o_3897),
  .I0(mux_o_3856),
  .I1(mux_o_3857),
  .S0(rad[5])
);
MUX2 mux_inst_3898 (
  .O(mux_o_3898),
  .I0(mux_o_3858),
  .I1(mux_o_3859),
  .S0(rad[5])
);
MUX2 mux_inst_3899 (
  .O(mux_o_3899),
  .I0(mux_o_3860),
  .I1(mux_o_3861),
  .S0(rad[5])
);
MUX2 mux_inst_3900 (
  .O(mux_o_3900),
  .I0(mux_o_3862),
  .I1(mux_o_3863),
  .S0(rad[5])
);
MUX2 mux_inst_3901 (
  .O(mux_o_3901),
  .I0(mux_o_3864),
  .I1(mux_o_3865),
  .S0(rad[5])
);
MUX2 mux_inst_3902 (
  .O(mux_o_3902),
  .I0(mux_o_3866),
  .I1(mux_o_3867),
  .S0(rad[5])
);
MUX2 mux_inst_3903 (
  .O(mux_o_3903),
  .I0(mux_o_3868),
  .I1(mux_o_3869),
  .S0(rad[5])
);
MUX2 mux_inst_3904 (
  .O(mux_o_3904),
  .I0(mux_o_3870),
  .I1(mux_o_3871),
  .S0(rad[5])
);
MUX2 mux_inst_3905 (
  .O(mux_o_3905),
  .I0(mux_o_3872),
  .I1(mux_o_3873),
  .S0(rad[5])
);
MUX2 mux_inst_3906 (
  .O(mux_o_3906),
  .I0(mux_o_3874),
  .I1(mux_o_3875),
  .S0(rad[6])
);
MUX2 mux_inst_3907 (
  .O(mux_o_3907),
  .I0(mux_o_3876),
  .I1(mux_o_3877),
  .S0(rad[6])
);
MUX2 mux_inst_3908 (
  .O(mux_o_3908),
  .I0(mux_o_3878),
  .I1(mux_o_3879),
  .S0(rad[6])
);
MUX2 mux_inst_3909 (
  .O(mux_o_3909),
  .I0(mux_o_3880),
  .I1(mux_o_3881),
  .S0(rad[6])
);
MUX2 mux_inst_3910 (
  .O(mux_o_3910),
  .I0(mux_o_3882),
  .I1(mux_o_3883),
  .S0(rad[6])
);
MUX2 mux_inst_3911 (
  .O(mux_o_3911),
  .I0(mux_o_3884),
  .I1(mux_o_3885),
  .S0(rad[6])
);
MUX2 mux_inst_3912 (
  .O(mux_o_3912),
  .I0(mux_o_3886),
  .I1(mux_o_3887),
  .S0(rad[6])
);
MUX2 mux_inst_3913 (
  .O(mux_o_3913),
  .I0(mux_o_3888),
  .I1(mux_o_3889),
  .S0(rad[6])
);
MUX2 mux_inst_3914 (
  .O(mux_o_3914),
  .I0(mux_o_3890),
  .I1(mux_o_3891),
  .S0(rad[6])
);
MUX2 mux_inst_3915 (
  .O(mux_o_3915),
  .I0(mux_o_3892),
  .I1(mux_o_3893),
  .S0(rad[6])
);
MUX2 mux_inst_3916 (
  .O(mux_o_3916),
  .I0(mux_o_3894),
  .I1(mux_o_3895),
  .S0(rad[6])
);
MUX2 mux_inst_3917 (
  .O(mux_o_3917),
  .I0(mux_o_3896),
  .I1(mux_o_3897),
  .S0(rad[6])
);
MUX2 mux_inst_3918 (
  .O(mux_o_3918),
  .I0(mux_o_3898),
  .I1(mux_o_3899),
  .S0(rad[6])
);
MUX2 mux_inst_3919 (
  .O(mux_o_3919),
  .I0(mux_o_3900),
  .I1(mux_o_3901),
  .S0(rad[6])
);
MUX2 mux_inst_3920 (
  .O(mux_o_3920),
  .I0(mux_o_3902),
  .I1(mux_o_3903),
  .S0(rad[6])
);
MUX2 mux_inst_3921 (
  .O(mux_o_3921),
  .I0(mux_o_3904),
  .I1(mux_o_3905),
  .S0(rad[6])
);
MUX2 mux_inst_3922 (
  .O(mux_o_3922),
  .I0(mux_o_3906),
  .I1(mux_o_3907),
  .S0(rad[7])
);
MUX2 mux_inst_3923 (
  .O(mux_o_3923),
  .I0(mux_o_3908),
  .I1(mux_o_3909),
  .S0(rad[7])
);
MUX2 mux_inst_3924 (
  .O(mux_o_3924),
  .I0(mux_o_3910),
  .I1(mux_o_3911),
  .S0(rad[7])
);
MUX2 mux_inst_3925 (
  .O(mux_o_3925),
  .I0(mux_o_3912),
  .I1(mux_o_3913),
  .S0(rad[7])
);
MUX2 mux_inst_3926 (
  .O(mux_o_3926),
  .I0(mux_o_3914),
  .I1(mux_o_3915),
  .S0(rad[7])
);
MUX2 mux_inst_3927 (
  .O(mux_o_3927),
  .I0(mux_o_3916),
  .I1(mux_o_3917),
  .S0(rad[7])
);
MUX2 mux_inst_3928 (
  .O(mux_o_3928),
  .I0(mux_o_3918),
  .I1(mux_o_3919),
  .S0(rad[7])
);
MUX2 mux_inst_3929 (
  .O(mux_o_3929),
  .I0(mux_o_3920),
  .I1(mux_o_3921),
  .S0(rad[7])
);
MUX2 mux_inst_3930 (
  .O(mux_o_3930),
  .I0(mux_o_3922),
  .I1(mux_o_3923),
  .S0(rad[8])
);
MUX2 mux_inst_3931 (
  .O(mux_o_3931),
  .I0(mux_o_3924),
  .I1(mux_o_3925),
  .S0(rad[8])
);
MUX2 mux_inst_3932 (
  .O(mux_o_3932),
  .I0(mux_o_3926),
  .I1(mux_o_3927),
  .S0(rad[8])
);
MUX2 mux_inst_3933 (
  .O(mux_o_3933),
  .I0(mux_o_3928),
  .I1(mux_o_3929),
  .S0(rad[8])
);
MUX2 mux_inst_3934 (
  .O(mux_o_3934),
  .I0(mux_o_3930),
  .I1(mux_o_3931),
  .S0(rad[9])
);
MUX2 mux_inst_3935 (
  .O(mux_o_3935),
  .I0(mux_o_3932),
  .I1(mux_o_3933),
  .S0(rad[9])
);
MUX2 mux_inst_3936 (
  .O(dout[30]),
  .I0(mux_o_3934),
  .I1(mux_o_3935),
  .S0(rad[10])
);
MUX2 mux_inst_3937 (
  .O(mux_o_3937),
  .I0(ram16sdp_inst_7_dout[31]),
  .I1(ram16sdp_inst_15_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3938 (
  .O(mux_o_3938),
  .I0(ram16sdp_inst_23_dout[31]),
  .I1(ram16sdp_inst_31_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3939 (
  .O(mux_o_3939),
  .I0(ram16sdp_inst_39_dout[31]),
  .I1(ram16sdp_inst_47_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3940 (
  .O(mux_o_3940),
  .I0(ram16sdp_inst_55_dout[31]),
  .I1(ram16sdp_inst_63_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3941 (
  .O(mux_o_3941),
  .I0(ram16sdp_inst_71_dout[31]),
  .I1(ram16sdp_inst_79_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3942 (
  .O(mux_o_3942),
  .I0(ram16sdp_inst_87_dout[31]),
  .I1(ram16sdp_inst_95_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3943 (
  .O(mux_o_3943),
  .I0(ram16sdp_inst_103_dout[31]),
  .I1(ram16sdp_inst_111_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3944 (
  .O(mux_o_3944),
  .I0(ram16sdp_inst_119_dout[31]),
  .I1(ram16sdp_inst_127_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3945 (
  .O(mux_o_3945),
  .I0(ram16sdp_inst_135_dout[31]),
  .I1(ram16sdp_inst_143_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3946 (
  .O(mux_o_3946),
  .I0(ram16sdp_inst_151_dout[31]),
  .I1(ram16sdp_inst_159_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3947 (
  .O(mux_o_3947),
  .I0(ram16sdp_inst_167_dout[31]),
  .I1(ram16sdp_inst_175_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3948 (
  .O(mux_o_3948),
  .I0(ram16sdp_inst_183_dout[31]),
  .I1(ram16sdp_inst_191_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3949 (
  .O(mux_o_3949),
  .I0(ram16sdp_inst_199_dout[31]),
  .I1(ram16sdp_inst_207_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3950 (
  .O(mux_o_3950),
  .I0(ram16sdp_inst_215_dout[31]),
  .I1(ram16sdp_inst_223_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3951 (
  .O(mux_o_3951),
  .I0(ram16sdp_inst_231_dout[31]),
  .I1(ram16sdp_inst_239_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3952 (
  .O(mux_o_3952),
  .I0(ram16sdp_inst_247_dout[31]),
  .I1(ram16sdp_inst_255_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3953 (
  .O(mux_o_3953),
  .I0(ram16sdp_inst_263_dout[31]),
  .I1(ram16sdp_inst_271_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3954 (
  .O(mux_o_3954),
  .I0(ram16sdp_inst_279_dout[31]),
  .I1(ram16sdp_inst_287_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3955 (
  .O(mux_o_3955),
  .I0(ram16sdp_inst_295_dout[31]),
  .I1(ram16sdp_inst_303_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3956 (
  .O(mux_o_3956),
  .I0(ram16sdp_inst_311_dout[31]),
  .I1(ram16sdp_inst_319_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3957 (
  .O(mux_o_3957),
  .I0(ram16sdp_inst_327_dout[31]),
  .I1(ram16sdp_inst_335_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3958 (
  .O(mux_o_3958),
  .I0(ram16sdp_inst_343_dout[31]),
  .I1(ram16sdp_inst_351_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3959 (
  .O(mux_o_3959),
  .I0(ram16sdp_inst_359_dout[31]),
  .I1(ram16sdp_inst_367_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3960 (
  .O(mux_o_3960),
  .I0(ram16sdp_inst_375_dout[31]),
  .I1(ram16sdp_inst_383_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3961 (
  .O(mux_o_3961),
  .I0(ram16sdp_inst_391_dout[31]),
  .I1(ram16sdp_inst_399_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3962 (
  .O(mux_o_3962),
  .I0(ram16sdp_inst_407_dout[31]),
  .I1(ram16sdp_inst_415_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3963 (
  .O(mux_o_3963),
  .I0(ram16sdp_inst_423_dout[31]),
  .I1(ram16sdp_inst_431_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3964 (
  .O(mux_o_3964),
  .I0(ram16sdp_inst_439_dout[31]),
  .I1(ram16sdp_inst_447_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3965 (
  .O(mux_o_3965),
  .I0(ram16sdp_inst_455_dout[31]),
  .I1(ram16sdp_inst_463_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3966 (
  .O(mux_o_3966),
  .I0(ram16sdp_inst_471_dout[31]),
  .I1(ram16sdp_inst_479_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3967 (
  .O(mux_o_3967),
  .I0(ram16sdp_inst_487_dout[31]),
  .I1(ram16sdp_inst_495_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3968 (
  .O(mux_o_3968),
  .I0(ram16sdp_inst_503_dout[31]),
  .I1(ram16sdp_inst_511_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3969 (
  .O(mux_o_3969),
  .I0(ram16sdp_inst_519_dout[31]),
  .I1(ram16sdp_inst_527_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3970 (
  .O(mux_o_3970),
  .I0(ram16sdp_inst_535_dout[31]),
  .I1(ram16sdp_inst_543_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3971 (
  .O(mux_o_3971),
  .I0(ram16sdp_inst_551_dout[31]),
  .I1(ram16sdp_inst_559_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3972 (
  .O(mux_o_3972),
  .I0(ram16sdp_inst_567_dout[31]),
  .I1(ram16sdp_inst_575_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3973 (
  .O(mux_o_3973),
  .I0(ram16sdp_inst_583_dout[31]),
  .I1(ram16sdp_inst_591_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3974 (
  .O(mux_o_3974),
  .I0(ram16sdp_inst_599_dout[31]),
  .I1(ram16sdp_inst_607_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3975 (
  .O(mux_o_3975),
  .I0(ram16sdp_inst_615_dout[31]),
  .I1(ram16sdp_inst_623_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3976 (
  .O(mux_o_3976),
  .I0(ram16sdp_inst_631_dout[31]),
  .I1(ram16sdp_inst_639_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3977 (
  .O(mux_o_3977),
  .I0(ram16sdp_inst_647_dout[31]),
  .I1(ram16sdp_inst_655_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3978 (
  .O(mux_o_3978),
  .I0(ram16sdp_inst_663_dout[31]),
  .I1(ram16sdp_inst_671_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3979 (
  .O(mux_o_3979),
  .I0(ram16sdp_inst_679_dout[31]),
  .I1(ram16sdp_inst_687_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3980 (
  .O(mux_o_3980),
  .I0(ram16sdp_inst_695_dout[31]),
  .I1(ram16sdp_inst_703_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3981 (
  .O(mux_o_3981),
  .I0(ram16sdp_inst_711_dout[31]),
  .I1(ram16sdp_inst_719_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3982 (
  .O(mux_o_3982),
  .I0(ram16sdp_inst_727_dout[31]),
  .I1(ram16sdp_inst_735_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3983 (
  .O(mux_o_3983),
  .I0(ram16sdp_inst_743_dout[31]),
  .I1(ram16sdp_inst_751_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3984 (
  .O(mux_o_3984),
  .I0(ram16sdp_inst_759_dout[31]),
  .I1(ram16sdp_inst_767_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3985 (
  .O(mux_o_3985),
  .I0(ram16sdp_inst_775_dout[31]),
  .I1(ram16sdp_inst_783_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3986 (
  .O(mux_o_3986),
  .I0(ram16sdp_inst_791_dout[31]),
  .I1(ram16sdp_inst_799_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3987 (
  .O(mux_o_3987),
  .I0(ram16sdp_inst_807_dout[31]),
  .I1(ram16sdp_inst_815_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3988 (
  .O(mux_o_3988),
  .I0(ram16sdp_inst_823_dout[31]),
  .I1(ram16sdp_inst_831_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3989 (
  .O(mux_o_3989),
  .I0(ram16sdp_inst_839_dout[31]),
  .I1(ram16sdp_inst_847_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3990 (
  .O(mux_o_3990),
  .I0(ram16sdp_inst_855_dout[31]),
  .I1(ram16sdp_inst_863_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3991 (
  .O(mux_o_3991),
  .I0(ram16sdp_inst_871_dout[31]),
  .I1(ram16sdp_inst_879_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3992 (
  .O(mux_o_3992),
  .I0(ram16sdp_inst_887_dout[31]),
  .I1(ram16sdp_inst_895_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3993 (
  .O(mux_o_3993),
  .I0(ram16sdp_inst_903_dout[31]),
  .I1(ram16sdp_inst_911_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3994 (
  .O(mux_o_3994),
  .I0(ram16sdp_inst_919_dout[31]),
  .I1(ram16sdp_inst_927_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3995 (
  .O(mux_o_3995),
  .I0(ram16sdp_inst_935_dout[31]),
  .I1(ram16sdp_inst_943_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3996 (
  .O(mux_o_3996),
  .I0(ram16sdp_inst_951_dout[31]),
  .I1(ram16sdp_inst_959_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3997 (
  .O(mux_o_3997),
  .I0(ram16sdp_inst_967_dout[31]),
  .I1(ram16sdp_inst_975_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3998 (
  .O(mux_o_3998),
  .I0(ram16sdp_inst_983_dout[31]),
  .I1(ram16sdp_inst_991_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_3999 (
  .O(mux_o_3999),
  .I0(ram16sdp_inst_999_dout[31]),
  .I1(ram16sdp_inst_1007_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_4000 (
  .O(mux_o_4000),
  .I0(ram16sdp_inst_1015_dout[31]),
  .I1(ram16sdp_inst_1023_dout[31]),
  .S0(rad[4])
);
MUX2 mux_inst_4001 (
  .O(mux_o_4001),
  .I0(mux_o_3937),
  .I1(mux_o_3938),
  .S0(rad[5])
);
MUX2 mux_inst_4002 (
  .O(mux_o_4002),
  .I0(mux_o_3939),
  .I1(mux_o_3940),
  .S0(rad[5])
);
MUX2 mux_inst_4003 (
  .O(mux_o_4003),
  .I0(mux_o_3941),
  .I1(mux_o_3942),
  .S0(rad[5])
);
MUX2 mux_inst_4004 (
  .O(mux_o_4004),
  .I0(mux_o_3943),
  .I1(mux_o_3944),
  .S0(rad[5])
);
MUX2 mux_inst_4005 (
  .O(mux_o_4005),
  .I0(mux_o_3945),
  .I1(mux_o_3946),
  .S0(rad[5])
);
MUX2 mux_inst_4006 (
  .O(mux_o_4006),
  .I0(mux_o_3947),
  .I1(mux_o_3948),
  .S0(rad[5])
);
MUX2 mux_inst_4007 (
  .O(mux_o_4007),
  .I0(mux_o_3949),
  .I1(mux_o_3950),
  .S0(rad[5])
);
MUX2 mux_inst_4008 (
  .O(mux_o_4008),
  .I0(mux_o_3951),
  .I1(mux_o_3952),
  .S0(rad[5])
);
MUX2 mux_inst_4009 (
  .O(mux_o_4009),
  .I0(mux_o_3953),
  .I1(mux_o_3954),
  .S0(rad[5])
);
MUX2 mux_inst_4010 (
  .O(mux_o_4010),
  .I0(mux_o_3955),
  .I1(mux_o_3956),
  .S0(rad[5])
);
MUX2 mux_inst_4011 (
  .O(mux_o_4011),
  .I0(mux_o_3957),
  .I1(mux_o_3958),
  .S0(rad[5])
);
MUX2 mux_inst_4012 (
  .O(mux_o_4012),
  .I0(mux_o_3959),
  .I1(mux_o_3960),
  .S0(rad[5])
);
MUX2 mux_inst_4013 (
  .O(mux_o_4013),
  .I0(mux_o_3961),
  .I1(mux_o_3962),
  .S0(rad[5])
);
MUX2 mux_inst_4014 (
  .O(mux_o_4014),
  .I0(mux_o_3963),
  .I1(mux_o_3964),
  .S0(rad[5])
);
MUX2 mux_inst_4015 (
  .O(mux_o_4015),
  .I0(mux_o_3965),
  .I1(mux_o_3966),
  .S0(rad[5])
);
MUX2 mux_inst_4016 (
  .O(mux_o_4016),
  .I0(mux_o_3967),
  .I1(mux_o_3968),
  .S0(rad[5])
);
MUX2 mux_inst_4017 (
  .O(mux_o_4017),
  .I0(mux_o_3969),
  .I1(mux_o_3970),
  .S0(rad[5])
);
MUX2 mux_inst_4018 (
  .O(mux_o_4018),
  .I0(mux_o_3971),
  .I1(mux_o_3972),
  .S0(rad[5])
);
MUX2 mux_inst_4019 (
  .O(mux_o_4019),
  .I0(mux_o_3973),
  .I1(mux_o_3974),
  .S0(rad[5])
);
MUX2 mux_inst_4020 (
  .O(mux_o_4020),
  .I0(mux_o_3975),
  .I1(mux_o_3976),
  .S0(rad[5])
);
MUX2 mux_inst_4021 (
  .O(mux_o_4021),
  .I0(mux_o_3977),
  .I1(mux_o_3978),
  .S0(rad[5])
);
MUX2 mux_inst_4022 (
  .O(mux_o_4022),
  .I0(mux_o_3979),
  .I1(mux_o_3980),
  .S0(rad[5])
);
MUX2 mux_inst_4023 (
  .O(mux_o_4023),
  .I0(mux_o_3981),
  .I1(mux_o_3982),
  .S0(rad[5])
);
MUX2 mux_inst_4024 (
  .O(mux_o_4024),
  .I0(mux_o_3983),
  .I1(mux_o_3984),
  .S0(rad[5])
);
MUX2 mux_inst_4025 (
  .O(mux_o_4025),
  .I0(mux_o_3985),
  .I1(mux_o_3986),
  .S0(rad[5])
);
MUX2 mux_inst_4026 (
  .O(mux_o_4026),
  .I0(mux_o_3987),
  .I1(mux_o_3988),
  .S0(rad[5])
);
MUX2 mux_inst_4027 (
  .O(mux_o_4027),
  .I0(mux_o_3989),
  .I1(mux_o_3990),
  .S0(rad[5])
);
MUX2 mux_inst_4028 (
  .O(mux_o_4028),
  .I0(mux_o_3991),
  .I1(mux_o_3992),
  .S0(rad[5])
);
MUX2 mux_inst_4029 (
  .O(mux_o_4029),
  .I0(mux_o_3993),
  .I1(mux_o_3994),
  .S0(rad[5])
);
MUX2 mux_inst_4030 (
  .O(mux_o_4030),
  .I0(mux_o_3995),
  .I1(mux_o_3996),
  .S0(rad[5])
);
MUX2 mux_inst_4031 (
  .O(mux_o_4031),
  .I0(mux_o_3997),
  .I1(mux_o_3998),
  .S0(rad[5])
);
MUX2 mux_inst_4032 (
  .O(mux_o_4032),
  .I0(mux_o_3999),
  .I1(mux_o_4000),
  .S0(rad[5])
);
MUX2 mux_inst_4033 (
  .O(mux_o_4033),
  .I0(mux_o_4001),
  .I1(mux_o_4002),
  .S0(rad[6])
);
MUX2 mux_inst_4034 (
  .O(mux_o_4034),
  .I0(mux_o_4003),
  .I1(mux_o_4004),
  .S0(rad[6])
);
MUX2 mux_inst_4035 (
  .O(mux_o_4035),
  .I0(mux_o_4005),
  .I1(mux_o_4006),
  .S0(rad[6])
);
MUX2 mux_inst_4036 (
  .O(mux_o_4036),
  .I0(mux_o_4007),
  .I1(mux_o_4008),
  .S0(rad[6])
);
MUX2 mux_inst_4037 (
  .O(mux_o_4037),
  .I0(mux_o_4009),
  .I1(mux_o_4010),
  .S0(rad[6])
);
MUX2 mux_inst_4038 (
  .O(mux_o_4038),
  .I0(mux_o_4011),
  .I1(mux_o_4012),
  .S0(rad[6])
);
MUX2 mux_inst_4039 (
  .O(mux_o_4039),
  .I0(mux_o_4013),
  .I1(mux_o_4014),
  .S0(rad[6])
);
MUX2 mux_inst_4040 (
  .O(mux_o_4040),
  .I0(mux_o_4015),
  .I1(mux_o_4016),
  .S0(rad[6])
);
MUX2 mux_inst_4041 (
  .O(mux_o_4041),
  .I0(mux_o_4017),
  .I1(mux_o_4018),
  .S0(rad[6])
);
MUX2 mux_inst_4042 (
  .O(mux_o_4042),
  .I0(mux_o_4019),
  .I1(mux_o_4020),
  .S0(rad[6])
);
MUX2 mux_inst_4043 (
  .O(mux_o_4043),
  .I0(mux_o_4021),
  .I1(mux_o_4022),
  .S0(rad[6])
);
MUX2 mux_inst_4044 (
  .O(mux_o_4044),
  .I0(mux_o_4023),
  .I1(mux_o_4024),
  .S0(rad[6])
);
MUX2 mux_inst_4045 (
  .O(mux_o_4045),
  .I0(mux_o_4025),
  .I1(mux_o_4026),
  .S0(rad[6])
);
MUX2 mux_inst_4046 (
  .O(mux_o_4046),
  .I0(mux_o_4027),
  .I1(mux_o_4028),
  .S0(rad[6])
);
MUX2 mux_inst_4047 (
  .O(mux_o_4047),
  .I0(mux_o_4029),
  .I1(mux_o_4030),
  .S0(rad[6])
);
MUX2 mux_inst_4048 (
  .O(mux_o_4048),
  .I0(mux_o_4031),
  .I1(mux_o_4032),
  .S0(rad[6])
);
MUX2 mux_inst_4049 (
  .O(mux_o_4049),
  .I0(mux_o_4033),
  .I1(mux_o_4034),
  .S0(rad[7])
);
MUX2 mux_inst_4050 (
  .O(mux_o_4050),
  .I0(mux_o_4035),
  .I1(mux_o_4036),
  .S0(rad[7])
);
MUX2 mux_inst_4051 (
  .O(mux_o_4051),
  .I0(mux_o_4037),
  .I1(mux_o_4038),
  .S0(rad[7])
);
MUX2 mux_inst_4052 (
  .O(mux_o_4052),
  .I0(mux_o_4039),
  .I1(mux_o_4040),
  .S0(rad[7])
);
MUX2 mux_inst_4053 (
  .O(mux_o_4053),
  .I0(mux_o_4041),
  .I1(mux_o_4042),
  .S0(rad[7])
);
MUX2 mux_inst_4054 (
  .O(mux_o_4054),
  .I0(mux_o_4043),
  .I1(mux_o_4044),
  .S0(rad[7])
);
MUX2 mux_inst_4055 (
  .O(mux_o_4055),
  .I0(mux_o_4045),
  .I1(mux_o_4046),
  .S0(rad[7])
);
MUX2 mux_inst_4056 (
  .O(mux_o_4056),
  .I0(mux_o_4047),
  .I1(mux_o_4048),
  .S0(rad[7])
);
MUX2 mux_inst_4057 (
  .O(mux_o_4057),
  .I0(mux_o_4049),
  .I1(mux_o_4050),
  .S0(rad[8])
);
MUX2 mux_inst_4058 (
  .O(mux_o_4058),
  .I0(mux_o_4051),
  .I1(mux_o_4052),
  .S0(rad[8])
);
MUX2 mux_inst_4059 (
  .O(mux_o_4059),
  .I0(mux_o_4053),
  .I1(mux_o_4054),
  .S0(rad[8])
);
MUX2 mux_inst_4060 (
  .O(mux_o_4060),
  .I0(mux_o_4055),
  .I1(mux_o_4056),
  .S0(rad[8])
);
MUX2 mux_inst_4061 (
  .O(mux_o_4061),
  .I0(mux_o_4057),
  .I1(mux_o_4058),
  .S0(rad[9])
);
MUX2 mux_inst_4062 (
  .O(mux_o_4062),
  .I0(mux_o_4059),
  .I1(mux_o_4060),
  .S0(rad[9])
);
MUX2 mux_inst_4063 (
  .O(dout[31]),
  .I0(mux_o_4061),
  .I1(mux_o_4062),
  .S0(rad[10])
);
endmodule //gowin_data_ram
