//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.01 (64-bit)
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Tue Mar 26 21:31:04 2024

module Gowin_SP_Instr (dout, clk, oce, ce, reset, wre, ad, din);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [13:0] ad;
input [31:0] din;

wire lut_f_0;
wire lut_f_1;
wire [26:0] spx9_inst_0_dout_w;
wire [8:0] spx9_inst_0_dout;
wire [26:0] spx9_inst_1_dout_w;
wire [8:0] spx9_inst_1_dout;
wire [26:0] spx9_inst_2_dout_w;
wire [8:0] spx9_inst_2_dout;
wire [26:0] spx9_inst_3_dout_w;
wire [8:0] spx9_inst_3_dout;
wire [26:0] spx9_inst_4_dout_w;
wire [17:9] spx9_inst_4_dout;
wire [26:0] spx9_inst_5_dout_w;
wire [17:9] spx9_inst_5_dout;
wire [26:0] spx9_inst_6_dout_w;
wire [17:9] spx9_inst_6_dout;
wire [26:0] spx9_inst_7_dout_w;
wire [17:9] spx9_inst_7_dout;
wire [29:0] sp_inst_8_dout_w;
wire [19:18] sp_inst_8_dout;
wire [29:0] sp_inst_9_dout_w;
wire [21:20] sp_inst_9_dout;
wire [29:0] sp_inst_10_dout_w;
wire [23:22] sp_inst_10_dout;
wire [29:0] sp_inst_11_dout_w;
wire [25:24] sp_inst_11_dout;
wire [29:0] sp_inst_12_dout_w;
wire [27:26] sp_inst_12_dout;
wire [29:0] sp_inst_13_dout_w;
wire [29:28] sp_inst_13_dout;
wire [29:0] sp_inst_14_dout_w;
wire [31:30] sp_inst_14_dout;
wire [15:0] sp_inst_15_dout_w;
wire [15:0] sp_inst_15_dout;
wire [15:0] sp_inst_16_dout_w;
wire [31:16] sp_inst_16_dout;
wire [31:0] sp_inst_17_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_14;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_31;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_48;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_65;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_82;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_99;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_116;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_133;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_150;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_167;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_184;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_201;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_218;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_235;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_252;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_269;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_286;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_303;
wire mux_o_310;
wire mux_o_320;
wire mux_o_330;
wire mux_o_340;
wire mux_o_350;
wire mux_o_360;
wire mux_o_370;
wire mux_o_380;
wire mux_o_390;
wire mux_o_400;
wire mux_o_410;
wire mux_o_420;
wire mux_o_430;
wire mux_o_440;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_0.INIT = 16'h0100;
LUT5 lut_inst_1 (
  .F(lut_f_1),
  .I0(ad[9]),
  .I1(ad[10]),
  .I2(ad[11]),
  .I3(ad[12]),
  .I4(ad[13])
);
defparam lut_inst_1.INIT = 32'h00040000;
SPX9 spx9_inst_0 (
    .DO({spx9_inst_0_dout_w[26:0],spx9_inst_0_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_0.READ_MODE = 1'b0;
defparam spx9_inst_0.WRITE_MODE = 2'b01;
defparam spx9_inst_0.BIT_WIDTH = 9;
defparam spx9_inst_0.BLK_SEL = 3'b000;
defparam spx9_inst_0.RESET_MODE = "SYNC";
defparam spx9_inst_0.INIT_RAM_00 = 288'hC67B3198C160B0182C166B31980D66B41B8C0673F1DEF17E3059AD07E401FF0F7CBC000D;
defparam spx9_inst_0.INIT_RAM_01 = 288'h0000000000000000000000000000000000000000000001000040003188F000C16630D82C;
defparam spx9_inst_0.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_20 = 288'hD0637418DD0637418DD063418A350AAD54A95429D4CA5522D166B258AC15EAE56AB0AA35;
defparam spx9_inst_0.INIT_RAM_21 = 288'h52A9168B3592C560AF572B5585500003418D000000000000000000000000000D0637418D;
defparam spx9_inst_0.INIT_RAM_22 = 288'hFF813218CC62B38085078381AC603184C620C20323F0884020001551A8556AA54AA14EA6;
defparam spx9_inst_0.INIT_RAM_23 = 288'h582BD5CAD561546A208FC221008FFCA5D8078FC221008C04B1122031987FE04FFF3BDFAD;
defparam spx9_inst_0.INIT_RAM_24 = 288'hC66B01A00CA85558B65128D42AB552A550A75329548BF5F2F578BB5D2E570B75A2CD64B1;
defparam spx9_inst_0.INIT_RAM_25 = 288'h552A550A75329548BF5F2F578BB5D2E570B75A2CD64B1582BD5CAD56157FE8402003599F;
defparam spx9_inst_0.INIT_RAM_26 = 288'h6660319AC6633400C06663198C06030198C656310EC7631880198C060B16AB65128D42AB;
defparam spx9_inst_0.INIT_RAM_27 = 288'h3B18C40633B0031ACD6663418CD6663198CCD633758CC66B3358CD0633199AC66035998C;
defparam spx9_inst_0.INIT_RAM_28 = 288'hC6EB75BCC663381A006067F198CC603001AC66B31998C666375A0CD6B319A00603158876;
defparam spx9_inst_0.INIT_RAM_29 = 288'h6031588763B18C40633B0031BADD6F319D8C660373F8CC66301800C6B331B8C6633318CC;
defparam spx9_inst_0.INIT_RAM_2A = 288'h066B598CDC6EB75BCC663381B9FC6633180C00001818D06335998C666375A0CD6B319A00;
defparam spx9_inst_0.INIT_RAM_2B = 288'h006B19ACC66631998DD6EB798CC670373F8CC66301800006B19ACC6663198CCC63331BAD;
defparam spx9_inst_0.INIT_RAM_2C = 288'h06637180C3B1D8C620319D8018DD6F341A0CC7630198DD6EB4198DC6030EC7631880C676;
defparam spx9_inst_0.INIT_RAM_2D = 288'h319D8C384667FFFF8402B33FECC06300EC763098C40633B0031BADD68331B8C066375BAD;
defparam spx9_inst_0.INIT_RAM_2E = 288'h3B18401FFFFE100ACCFFFFD980C601D8EC6131880C676308033F8C467FC00763B184C620;
defparam spx9_inst_0.INIT_RAM_2F = 288'h3B1D8C2631018CEC61C263199FFFFE100ACCFFE100ACCFFB0180C066030EC763098C4063;
defparam spx9_inst_0.INIT_RAM_30 = 288'h1018CEC61007FFFFFFC201599FFFFB3318CC6663198CCC6331998C6633318CC6603180C4;
defparam spx9_inst_0.INIT_RAM_31 = 288'h62FFF0805667FFFECCC6331998C6633318CC6663198CCC6331980C603198AC43B1D8C263;
defparam spx9_inst_0.INIT_RAM_32 = 288'h6633318CC6663198CCC6331998C6633018C06331588763B184C620319D8C200FFFFFFEC4;
defparam spx9_inst_0.INIT_RAM_33 = 288'h31880C676308000004C2B31988C3B1D8C2631018CEC61007FFFEC462FFF0805667FD998C;
defparam spx9_inst_0.INIT_RAM_34 = 288'h66EB39ACE66F300F80D73359800603319800FF811980C6660199806631D8CC5621D8EC61;
defparam spx9_inst_0.INIT_RAM_35 = 288'h06335980C0063358CDC63331ACC6680199CCC673B5ACE66B333ECC6663198CC03E8398CE;
defparam spx9_inst_0.INIT_RAM_36 = 288'hD60319A00621D8EC6131880C67630E10180C6633318CCFFE13198CC6330018CC6631998D;
defparam spx9_inst_0.INIT_RAM_37 = 288'h6632D94C96431D8CC5621D8EC6131880C67630E10199F6633318CC6663199FFC2333FE04;
defparam spx9_inst_0.INIT_RAM_38 = 288'hC6333018CD6631998DD6037198CD633718CC66033580C66B3319AC66B3000C066331998C;
defparam spx9_inst_0.INIT_RAM_39 = 288'h6633318CCFFE118A0603E3198006663198CCC6333FF84C663198006663198CCC6333FF84;
defparam spx9_inst_0.INIT_RAM_3A = 288'h66001998C6633318CCFFE118A0603E3198006663198CCC6333FF84628180F8C66001998C;
defparam spx9_inst_0.INIT_RAM_3B = 288'h6663199FF02001998C6633318CCFFE118A0603E3198006663198CCC6333FF84628180F8C;
defparam spx9_inst_0.INIT_RAM_3C = 288'hC6EB19B8C66634198DD633718CC6663198CCD663319CC6763199AD0633400C0666319800;
defparam spx9_inst_0.INIT_RAM_3D = 288'h0663758CDC63331A0CC6EB19B8C6633318CC666B3198CE633B18CCD68319A00607FF1A0C;
defparam spx9_inst_0.INIT_RAM_3E = 288'h621D8EC631018CEC61C20333F8CD633598CCC6333FF84667FC09AC063340000FF813FF8D;
defparam spx9_inst_0.INIT_RAM_3F = 288'h06B3300CCC6B331B8CC66319980666341ACCC6835998D66637580CC6E31998D06B3180C0;

SPX9 spx9_inst_1 (
    .DO({spx9_inst_1_dout_w[26:0],spx9_inst_1_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_1.READ_MODE = 1'b0;
defparam spx9_inst_1.WRITE_MODE = 2'b01;
defparam spx9_inst_1.BIT_WIDTH = 9;
defparam spx9_inst_1.BLK_SEL = 3'b001;
defparam spx9_inst_1.RESET_MODE = "SYNC";
defparam spx9_inst_1.INIT_RAM_00 = 288'hC0030EC7631880C676006359ACCCFE33198C6600198AC621D8EC631018CEC0066631998D;
defparam spx9_inst_1.INIT_RAM_01 = 288'h3B18C40633B000580C3B1D8C620319D800203B1D8C620319D8018C061D8EC631018CEC00;
defparam spx9_inst_1.INIT_RAM_02 = 288'h66E3018CCD6337598CF6637180C6033318CCC033188763B18C40633B00059AC063358876;
defparam spx9_inst_1.INIT_RAM_03 = 288'h00333198CC6031988C3B1D8C620319D8018DE6837180CC76301800C6EB7180CC6E30198D;
defparam spx9_inst_1.INIT_RAM_04 = 288'h6663198CCC6333FF84667FC09AC0633400C43B1D8C2631018CEC00C6B3419AC0663718CC;
defparam spx9_inst_1.INIT_RAM_05 = 288'h66B3000C06633001FF0233018CCC033300CC63B198AC43B1D8C2631018CEC61C20333ECC;
defparam spx9_inst_1.INIT_RAM_06 = 288'h6663598CD00333998CE76B59CCD6667D98CCC63319807D07319CCDD67359CCDE601F01AE;
defparam spx9_inst_1.INIT_RAM_07 = 288'h1018CEC61C203018CC6663199FFC2633198C66003198CC63331A0C66B301800C66B19B8C;
defparam spx9_inst_1.INIT_RAM_08 = 288'h66E3198CC066B018CD6663358CD6600180CC6633318CC65B2992C863B198AC43B1D8C263;
defparam spx9_inst_1.INIT_RAM_09 = 288'hC6331998C667FF098CC633000CCC6331998C667FF098C6660319ACC63331BAC06E3319AC;
defparam spx9_inst_1.INIT_RAM_0A = 288'hC633000CCC6331998C667FF08C50301F18CC0033318CC6663199FFC23140C07C633000CC;
defparam spx9_inst_1.INIT_RAM_0B = 288'hC23140C07C633000CCC6331998C667FF08C50301F18CC0033318CC6663199FFC23140C07;
defparam spx9_inst_1.INIT_RAM_0C = 288'hC633199ACC663398CEC63335A0C6680180CCC633000CCC6333FE040033318CC6663199FF;
defparam spx9_inst_1.INIT_RAM_0D = 288'h6663198CCD663319CC6763199AD0633400C0FFE34198DD633718CCC68331BAC66E3198CC;
defparam spx9_inst_1.INIT_RAM_0E = 288'hE60359D80667FF08CCFF813580C6680001FF027FF1A0CC6EB19B8C66634198DD633718CC;
defparam spx9_inst_1.INIT_RAM_0F = 288'h3B1D8C620319D8C3840667F19AC66B31998C6667D9B8D66000000000001998C566000FA0;
defparam spx9_inst_1.INIT_RAM_10 = 288'h66310EC763098C40633B003180C3B1D8C620319D80180061D8EC631018CED846633018C0;
defparam spx9_inst_1.INIT_RAM_11 = 288'h006B318CCC6B33598C66635998D66237FEC43B1D8C2631018CEC6100635988DFFE019980;
defparam spx9_inst_1.INIT_RAM_12 = 288'h66B13FF8466003FF84667FD80C060310EC763098C40633B18709ACC63335ACDC6331980C;
defparam spx9_inst_1.INIT_RAM_13 = 288'hC26B3182C66B10EC763098C40633B18401FFC263198C43B1D8C2631018CEC61007FF58CC;
defparam spx9_inst_1.INIT_RAM_14 = 288'hC06319B8D660018AC43B1D8C620319D8C200FFE13580C66B10EC763098C40633B18401FF;
defparam spx9_inst_1.INIT_RAM_15 = 288'h66633190C6030188763B18C40633B613598C6633318CCC6E3199ACC633B1CCCC6B30000C;
defparam spx9_inst_1.INIT_RAM_16 = 288'h66635998DC663318CCC6B331B8CC63331ACCC6E33198C66635998DC663318CC66633190C;
defparam spx9_inst_1.INIT_RAM_17 = 288'h666341ACCC0631998D0663598C43B1D8C620319D8018D66637198CC63331ACCC6E33198C;
defparam spx9_inst_1.INIT_RAM_18 = 288'h0663999ADC67B00F80E78331CCCC6F300F80D70331ACCC6836198D06B33018C66634198D;
defparam spx9_inst_1.INIT_RAM_19 = 288'hC663199ADC67B00F80E78331CCCC6E31998DC64331BED03E839E0DD7337598CF601F01CF;
defparam spx9_inst_1.INIT_RAM_1A = 288'h31880C67630803FEC4007FD8980663318A8C3B1D8C2631018CEC00C6837190CC6E3219AD;
defparam spx9_inst_1.INIT_RAM_1B = 288'h006375A0CC7731980EC6830018DD68331C0CE63301D8D0660198CC6663418CD62B10EC76;
defparam spx9_inst_1.INIT_RAM_1C = 288'h3B1D8C620319D8018DD68331DCC6603B1A0C006375A0CC703398CC0763419806633318CC;
defparam spx9_inst_1.INIT_RAM_1D = 288'hC6330018DD68331DCC6603B1A0C006375A0CC703398CC07634198066331998D063358AC4;
defparam spx9_inst_1.INIT_RAM_1E = 288'hC6030EC7631880C676006375A0CC7731980EC6830018DD68331C0CE63301D8D0660198CC;
defparam spx9_inst_1.INIT_RAM_1F = 288'hC60331D8C066379BADF6E30198EC6033018C663018AC43B1D8C620319D8018DD6EB4198D;
defparam spx9_inst_1.INIT_RAM_20 = 288'h66635998D666B718CCC6B331ACCD6E31998D660031ACCD683318CCC6B33018C666379A0D;
defparam spx9_inst_1.INIT_RAM_21 = 288'hC6B335B8C66635998D666B4198C666359800C6B335B8C6663599AC06635998D666B4198C;
defparam spx9_inst_1.INIT_RAM_22 = 288'h31880C67600601998D06B331A0D6660198C43B1D8C620319D8018D666B4198C666359800;
defparam spx9_inst_1.INIT_RAM_23 = 288'h319D8018DE6B34198E063331BAD5683188763B18C40633B0031ACCD6B331ACC62B10EC76;
defparam spx9_inst_1.INIT_RAM_24 = 288'h6601F41CC67635998D06B31998C163018AC43B1D8C2631018CEC00C6EB55A0C3B1D8C620;
defparam spx9_inst_1.INIT_RAM_25 = 288'h6660318CCC6B331BAC06637598C66637598C66635998D6663718CCC6B331ACC6663318CC;
defparam spx9_inst_1.INIT_RAM_26 = 288'hC03331A0D666341ACCC6835998DD6C3598C43B1D8C620319D8C200000131ACCC6B331A0D;
defparam spx9_inst_1.INIT_RAM_27 = 288'h31880C67600635998DD60331B8C660031ACCC6E33198C6660198C5621D8EC631018CEC00;
defparam spx9_inst_1.INIT_RAM_28 = 288'hC63331ACC003118CC5621D8EC6131880C676308031A0D066359ACC0031198AC621D8EC61;
defparam spx9_inst_1.INIT_RAM_29 = 288'h422930ACC6663199806600188CCD63319AAC621D8EC6131880C676308031ACCC6E3319AC;
defparam spx9_inst_1.INIT_RAM_2A = 288'hC633000CCC633188763B18C40633B184018D068331ACD667FD08A4C2B3199AC0633401FF;
defparam spx9_inst_1.INIT_RAM_2B = 288'h3B184C620319D8018D66637198CC6333018C6633318CC621D8EC631018CEC00CFE3198CC;
defparam spx9_inst_1.INIT_RAM_2C = 288'hC663019FF027FC098503333FE84526174CCD66333198CC663198CCC633199AC662B51876;
defparam spx9_inst_1.INIT_RAM_2D = 288'hFF8130ACCFFA110980C6633180CFF813FE04C2E3199FF422130ACC6663199FF42213018C;
defparam spx9_inst_1.INIT_RAM_2E = 288'hC663198CCC6331988C3B1D8C2631018CEC61007FC09FF02017FE8442603198CC6033FE04;
defparam spx9_inst_1.INIT_RAM_2F = 288'h6633318CCFFA110985667FD0884C0633198C067FC09FF026140CCCFFA11098566333198C;
defparam spx9_inst_1.INIT_RAM_30 = 288'h020140DFF42213018CC663019FF027FC098503333FE8442603198CC6033FE04FF8130B8C;
defparam spx9_inst_1.INIT_RAM_31 = 288'h006B018CD66633180C00333198C066341B8C061D8EC631018CEC61C2331998C067FC09FF;
defparam spx9_inst_1.INIT_RAM_32 = 288'h66E359B8C066379BADF6B3819AC06335998CC603000CCC663018C662B10EC7631880C676;
defparam spx9_inst_1.INIT_RAM_33 = 288'hE6633D98EC63335B8CC63331B8C66310EC7631880C676006341B8C060031A0DC6033580C;
defparam spx9_inst_1.INIT_RAM_34 = 288'hD6F30198EC63331B8C66310EC7631880C67600637188CD6E3318CCD6F33182CC763199AD;
defparam spx9_inst_1.INIT_RAM_35 = 288'hF663B18CCC6E3198C43B1D8C620319D8018DC62331BAD66EB3198CC63335BCC0663B18CC;
defparam spx9_inst_1.INIT_RAM_36 = 288'hC663199ADC663318CCD6E33198C666B7198CC63335B8CC663199ADE63B31D8C666B7998C;
defparam spx9_inst_1.INIT_RAM_37 = 288'h319D8018DE6837180CC76301800C6EB7180CC6E30198066310EC7631880C6760063519AD;
defparam spx9_inst_1.INIT_RAM_38 = 288'hC66B3188CC6E3198CC461D8EC631018CED84C6633198CD6631198DC6331988C3B1D8C620;
defparam spx9_inst_1.INIT_RAM_39 = 288'h31880C676006375A8CC6A30EC7631880C676006375A8CC6A30EC7631880C676C2633198C;
defparam spx9_inst_1.INIT_RAM_3A = 288'h3B18C40633B003598CF6EB51BAFD6B375DAD66E3319ACC62331B8C6633358CC56A30EC76;
defparam spx9_inst_1.INIT_RAM_3B = 288'h3B184C620319D801ACE67B75A8DD7EB59B8CC66B3188CC6E31998EC633199AC662B51876;
defparam spx9_inst_1.INIT_RAM_3C = 288'h66031980C66230EC763098C40633B184018D06335998C667FF09A566E319800603311876;
defparam spx9_inst_1.INIT_RAM_3D = 288'h66031980C6033018CC0633019FFC2331980C66031980C6033019FFC2331980C66031980C;
defparam spx9_inst_1.INIT_RAM_3E = 288'h467FF098C6600180763B184C620319D8C200FF813FF846667F198C46003FFFFC233180C0;
defparam spx9_inst_1.INIT_RAM_3F = 288'hC68319ACCC6333FE844261719AC66E319800607FD0884C68319ACCC63331BCC67631998D;

SPX9 spx9_inst_2 (
    .DO({spx9_inst_2_dout_w[26:0],spx9_inst_2_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_2.READ_MODE = 1'b0;
defparam spx9_inst_2.WRITE_MODE = 2'b01;
defparam spx9_inst_2.BIT_WIDTH = 9;
defparam spx9_inst_2.BLK_SEL = 3'b010;
defparam spx9_inst_2.RESET_MODE = "SYNC";
defparam spx9_inst_2.INIT_RAM_00 = 288'hC60331BAD66E301980C6033000C621D8EC631018CEC61007FD0884C2B31998CC6633188C;
defparam spx9_inst_2.INIT_RAM_01 = 288'h06635998E066379A0CC6B331C0CC6EB75A0CC6E301980C63331BCD06635998E066375ACD;
defparam spx9_inst_2.INIT_RAM_02 = 288'h666375A6D666375A2D666341ACCC6835998D06B331BAD16B3188763B18C40633B0031BCD;
defparam spx9_inst_2.INIT_RAM_03 = 288'hC033188763B18C40633B0031BAD066341800C6EB4198D0660198C43B1D8C620319D80180;
defparam spx9_inst_2.INIT_RAM_04 = 288'h3B18C40633B0031BADE6834198EC60331BAD066341800C6EB75A0CC6E30198DD68331A0C;
defparam spx9_inst_2.INIT_RAM_05 = 288'h06637198C066379ACD0663818C43B1D8C620319DB08CC60001980CC06B1998D063018876;
defparam spx9_inst_2.INIT_RAM_06 = 288'h621D8EC631018CEC61000010984C2B331A0DC6631988C3B1D8C2631018CEC00C6EB75B8C;
defparam spx9_inst_2.INIT_RAM_07 = 288'h6663718CCC6B331ACCC6E319980666B318CCC6B331ACCC6E31998D66E335ACDC633198AC;
defparam spx9_inst_2.INIT_RAM_08 = 288'h3B184C620319DB080062B10EC7631880C6760060199ACC63331ACCC6B331B8C66635998D;
defparam spx9_inst_2.INIT_RAM_09 = 288'h46B3318CCFFA1109C5C3633598C666B51B8E6600181FF4221001AC06337580C66B158876;
defparam spx9_inst_2.INIT_RAM_0A = 288'hC63335A8DC0233FEC4C2E33598C666B51A006033318CC0067D19FF422130B8CD663199AD;
defparam spx9_inst_2.INIT_RAM_0B = 288'h4261719ACC63335A8D666319800FFA1109C5F361F19ACC63335A8DC7EB318CCD6A371DAC;
defparam spx9_inst_2.INIT_RAM_0C = 288'h31880C67630E101800007FD0884007FD0884C0233FE844261719ACC63335A8DCFA33FE84;
defparam spx9_inst_2.INIT_RAM_0D = 288'h66000000000001998C567FD0884CFB371ACC0000000000033318ECC6837180CFF9D8EC61;
defparam spx9_inst_2.INIT_RAM_0E = 288'h6663159FF422100ACCC62333ECDC6B3000000000000CCC62B3FE8442315998C4667D9B8D;
defparam spx9_inst_2.INIT_RAM_0F = 288'h02FFC0805CFB371ACC0000000000033318ACFFA11098566330199F66E359800000000000;
defparam spx9_inst_2.INIT_RAM_10 = 288'h020173ECDC6B3000000000000CCC61B3FE0402E7D9B8D66000000000001998C367FFFE04;
defparam spx9_inst_2.INIT_RAM_11 = 288'h00613198C6600019FF422131A0C66E3418CD62B10EC763098C40633B61018763B18FFFFF;
defparam spx9_inst_2.INIT_RAM_12 = 288'hC2E3319AC66337FE844261758CC66E0318CC00301988C00613198C66001980CD60319AC4;
defparam spx9_inst_2.INIT_RAM_13 = 288'h00033FE844263418CDC68319AC5621D8EC6131880C67630E1019AC66335998C667FD0884;
defparam spx9_inst_2.INIT_RAM_14 = 288'h422130BAC6663718CCC06319800603311800C263318CC0033019AC063358800C263318CC;
defparam spx9_inst_2.INIT_RAM_15 = 288'hD60319AC5621D8EC6131880C67630E1019AC66335998C667FD0884C2E3358CCC6E3199FF;
defparam spx9_inst_2.INIT_RAM_16 = 288'h621D8EC6131880C67630E10198D66B31988C00613198C663100184C66319800067FD0884;
defparam spx9_inst_2.INIT_RAM_17 = 288'h3098C40633B187080CC6B3598C400613198C663100184C66319800067FD0884D60319AC5;
defparam spx9_inst_2.INIT_RAM_18 = 288'h0033018CC066B0198D66001980C66033580CC6E3199AC0663718CCD60331ACC60310EC76;
defparam spx9_inst_2.INIT_RAM_19 = 288'h6663358CCD6B319B8D063371A0C66803580C66EB018CDD60319ACCC66B198CD0033018C0;
defparam spx9_inst_2.INIT_RAM_1A = 288'hFFA1108006663358CCD6B319B8D063371A0C66801998CD63335ACC66E3418CDC68319A00;
defparam spx9_inst_2.INIT_RAM_1B = 288'h30E11999FC66B198CD666319800FFA1108006663358CCD6B319BAC66E31998D063340000;
defparam spx9_inst_2.INIT_RAM_1C = 288'h42193FEC4FFE13198C66313FF84C66319800067FD0864D60319AC5621D8EC6131880C676;
defparam spx9_inst_2.INIT_RAM_1D = 288'h32617198C467FD0864C2E3119FF42190EC763098C40633B187080CFFA10C9FF623140DFF;
defparam spx9_inst_2.INIT_RAM_1E = 288'h323174D87C6733188CC7631998DD6631198DC633000C0FFA10C9FF421930B8CC6233FE84;
defparam spx9_inst_2.INIT_RAM_1F = 288'hC2A33FF84C633000C0FFA10C9FF42190EC763098C40633B187080CC68319ACCC6333FE84;
defparam spx9_inst_2.INIT_RAM_20 = 288'h30E10198D06335998C667FD0864C2A33FF84C633000C0FFA10C98D06335998C667FD0864;
defparam spx9_inst_2.INIT_RAM_21 = 288'hC663199FF42190000CFFA10C9AC06337008CFFA10C985C663198C5621D8EC6131880C676;
defparam spx9_inst_2.INIT_RAM_22 = 288'h66003FFFFFFA10C980C66B3198CC63331B8C467FD0864C2E3318CC007FF08CC66233FF84;
defparam spx9_inst_2.INIT_RAM_23 = 288'h66B3318CCFFE134ACC6680181AC06335988CFFE13198C667FD0864C0233FE8432617198C;
defparam spx9_inst_2.INIT_RAM_24 = 288'h467FD0864C2E3318CC00033FE8432003FF84D2B319ACC467FF098CC6333580C668031A0C;
defparam spx9_inst_2.INIT_RAM_25 = 288'hFFE0319ACC663318CCC6E3119FF421930B8CC633001FFFFA10C980C66B3198CC63331B8C;
defparam spx9_inst_2.INIT_RAM_26 = 288'hFF813FE04C68319BFF421918AC43B1D8C2631018CEC61C2030000CFFA10C9FF4219001FF;
defparam spx9_inst_2.INIT_RAM_27 = 288'hC60B19ACCC6333FF8466313FF84C663198C4FFE13198C66313FF84C66319800067FD0864;
defparam spx9_inst_2.INIT_RAM_28 = 288'h42193FF8D06337FE84323158AC43B1D8C2631018CEC61C2033FF8466333598C1633599AC;
defparam spx9_inst_2.INIT_RAM_29 = 288'h421931A0C66B1588763B184C620319D8C384067FF09ACC66319AC4FFE13198C6600019FF;
defparam spx9_inst_2.INIT_RAM_2A = 288'h32317FEC4D60319A00FFA10C8C5FFB13580C66B13FF84C663198C4FFE13198C6600019FF;
defparam spx9_inst_2.INIT_RAM_2B = 288'hFFA10C8C562B10EC763098C40633B187080CFFA10C800FFA10C8C5FFB13580C66803FE84;
defparam spx9_inst_2.INIT_RAM_2C = 288'h66230EC763098C40633B187080CFFFFD88C4FFE13198C6600019FF42193FE04C68319BFF;
defparam spx9_inst_2.INIT_RAM_2D = 288'hC763F186CFFA10C8C5621D8EE763098C40633B187098C6600019FF421931A0C66E3418CD;
defparam spx9_inst_2.INIT_RAM_2E = 288'hC66319800067FD0864FFA10C9FF42193FE843260119FFC26959B8CC633198CD6733F198D;
defparam spx9_inst_2.INIT_RAM_2F = 288'hFFE13198C666DC188DFFE1318CC6663198CCC6330000CFFA10C9AC06337008CFFE134ACD;
defparam spx9_inst_2.INIT_RAM_30 = 288'hFFE13198C666DC188DFFE13198C66331D88CFFE13198C666DC188DFFE13198C66331D88C;
defparam spx9_inst_2.INIT_RAM_31 = 288'h467FF098CC63336E0C46FFF098CC633198EC467FF098CC63336E0C46FFF098C66331D88C;
defparam spx9_inst_2.INIT_RAM_32 = 288'h66EB018CDC03331A0C66E01998D0633598EC467FF098CC63336E0C46FFF098CC633198EC;
defparam spx9_inst_2.INIT_RAM_33 = 288'h6633318CC6663198CCC6330000CFFA10C9806633018000663418CDC68319B8D063371A0C;
defparam spx9_inst_2.INIT_RAM_34 = 288'hC6330000CFFA10C9AC06337008CFFE134ACDC66319800FF8130ACC6663198CCC6331998C;
defparam spx9_inst_2.INIT_RAM_35 = 288'hFFE13198C666DC188DFFE13198C66331D88CFFE13198C666DC188DFFE1318CC6663198CC;
defparam spx9_inst_2.INIT_RAM_36 = 288'h467FF098CC63336E0C46FFF098CC633198EC467FF098CC63336E0C46FFF098C66331D88C;
defparam spx9_inst_2.INIT_RAM_37 = 288'h66EB018CDC03331A0C66E01998D0633598EC467FF098CC63336E0C46FFF098CC633198EC;
defparam spx9_inst_2.INIT_RAM_38 = 288'h6633318CC6663198CCC6330000CFFA10C9806633018000663418CDC68319B8D063371A0C;
defparam spx9_inst_2.INIT_RAM_39 = 288'hC6733198C67637598C7633589FFC263318CCC0233FF84D2B37198C6600018CCC6331998C;
defparam spx9_inst_2.INIT_RAM_3A = 288'h6633198CC667FC0985667FD0864D60319A000633318CC666319800067FD0864C0633598C;
defparam spx9_inst_2.INIT_RAM_3B = 288'h62B10EC763098C40633B9D8C384067FD086462B198FFF421918AC663B3198CC6633198CC;
defparam spx9_inst_2.INIT_RAM_3C = 288'h621D8EC6131880C67630E1019FF62313FF84C66319800067FD0864FFE3418CDFFA10C8C5;
defparam spx9_inst_2.INIT_RAM_3D = 288'h667FD086400033FE84326B018CD62B10EC763098C40633B1870800FF8130ACCFFE1198C5;
defparam spx9_inst_2.INIT_RAM_3E = 288'h421930ACC66633598C6663718CC66233FF84C663198CC467FF098CC6331988CFFE13198C;
defparam spx9_inst_2.INIT_RAM_3F = 288'h6600019FF42193580C66B1588763B184C620319D8C384067FF09A566337FE843261599FF;

SPX9 spx9_inst_3 (
    .DO({spx9_inst_3_dout_w[26:0],spx9_inst_3_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_3.READ_MODE = 1'b0;
defparam spx9_inst_3.WRITE_MODE = 2'b01;
defparam spx9_inst_3.BIT_WIDTH = 9;
defparam spx9_inst_3.BLK_SEL = 3'b011;
defparam spx9_inst_3.RESET_MODE = "SYNC";
defparam spx9_inst_3.INIT_RAM_00 = 288'hC2B31988CFFE1198CCD6633198C66637598C76637198C66313FF84C663198C4FFE13198C;
defparam spx9_inst_3.INIT_RAM_01 = 288'h063371A0C66B13FF84C663198C4FFE13198C6631588763B184C620319D8C384067FD0864;
defparam spx9_inst_3.INIT_RAM_02 = 288'h0600019FF42193FE84327FD0864C0331988CFFE13198C6633018000663418CDC68319B8D;
defparam spx9_inst_3.INIT_RAM_03 = 288'hC6333FE843261719AC06335998CC60331BADC60331B8C066379ACDC60331CCC006361B8C;
defparam spx9_inst_3.INIT_RAM_04 = 288'h00033FE84326B018CD62B10EC763098C40633B187080CC6F375AEDC60331D8C0667D98CC;
defparam spx9_inst_3.INIT_RAM_05 = 288'hE6EB7DA0CC703001AC0633700CCD60319B8D063371BCD068331C0CC033189FFC263318CC;
defparam spx9_inst_3.INIT_RAM_06 = 288'h32000018DE6834198E066379BADF68331C0C006379A0D06638198DE6EB7DA0CC7030018D;
defparam spx9_inst_3.INIT_RAM_07 = 288'h660331A0DC60331A0DC60331A0DC6030EC763098C40633B187080CC6837180C00033FE84;
defparam spx9_inst_3.INIT_RAM_08 = 288'h66E3198CCC63331BAD66637580C6680198CCC683419FF42193FF8DE683419AEC67B19A00;
defparam spx9_inst_3.INIT_RAM_09 = 288'h667FD0844D6633980C6763598006633000CC066B018CD66631998DE683419AEC67B19B8D;
defparam spx9_inst_3.INIT_RAM_0A = 288'h00033FE84226B018CD62B10EC763098C40633B187080CD60319ACCC63331ACDC6331998C;
defparam spx9_inst_3.INIT_RAM_0B = 288'h3B184C620319D8C3840600019FF4211001FFC26B018CD007FE09AC0633589FFC263318CC;
defparam spx9_inst_3.INIT_RAM_0C = 288'hD60319AC5621D8EC6131880C67630E1001FF421130ACC66233FF8D068331A0D063158876;
defparam spx9_inst_3.INIT_RAM_0D = 288'h663371DAC066B598CD00301998C6600180CC067FD084460313FF84C66319800067FD0844;
defparam spx9_inst_3.INIT_RAM_0E = 288'h30E1019FF4211358CC66B3318CCFFE118A06D63319BFF421131A0C66B3318CCC6EB79BAC;
defparam spx9_inst_3.INIT_RAM_0F = 288'h6600180CC067FD084460313FF84C66319800067FD0844D60319AC5621D8EC6131880C676;
defparam spx9_inst_3.INIT_RAM_10 = 288'h066B598CDC763358CC66EB3198CE60339CCC6763758CC6680181FFC23140DAC66335998C;
defparam spx9_inst_3.INIT_RAM_11 = 288'h31880C67630E1019FF4211358CC66B3318CCFFA10898D06335998C66003FE84227170DAC;
defparam spx9_inst_3.INIT_RAM_12 = 288'h30E1019FFC26B018CDFFB13FE8422313FF84C66319800067FD0844D60319AC5621D8EC61;
defparam spx9_inst_3.INIT_RAM_13 = 288'hFFE13580C66FFD89FF421130ACC66233FF8D068331A0D0630180C5621D8EC6131880C676;
defparam spx9_inst_3.INIT_RAM_14 = 288'h663371A0C66B3318CCC6EB79BAC663371DAC066B598CD00301998C6600180CC067FD0844;
defparam spx9_inst_3.INIT_RAM_15 = 288'h6281B58CC66B3318CC00301980CFFA1089FF4211358CC66B3318CCFFA1089FFC23140DAC;
defparam spx9_inst_3.INIT_RAM_16 = 288'h007FD0844E2E1B580CD6B319B8EC66B198CDD663319CC0673998CEC6EB198CD00303FF84;
defparam spx9_inst_3.INIT_RAM_17 = 288'hC20300A063B1D8C2631018CEC61C2033FE84226B198CD6663199FF421131A0C66B3318CC;
defparam spx9_inst_3.INIT_RAM_18 = 288'h3B184C620319D8C384007FF080CC2B31980C66031980C6663019FFC2333FF84060140DFF;
defparam spx9_inst_3.INIT_RAM_19 = 288'h00303FE842231588763B184C620319DB080C6031588763B18C40633B187080CFFB158876;
defparam spx9_inst_3.INIT_RAM_1A = 288'h0633400C0D61319ACCC633359CCC6EB018CDC76B018CD00303584C66B3318CCC06B018CD;
defparam spx9_inst_3.INIT_RAM_1B = 288'h30E101980066B098CD6663199FF421118BC6C3E33580C66E3B580C66EB319CC0633B1BAC;
defparam spx9_inst_3.INIT_RAM_1C = 288'hFFA10880563118EC763098C40633B18401FFC20300BFF421100AC6231D8EC6131880C676;
defparam spx9_inst_3.INIT_RAM_1D = 288'h3B1D8C2631018CEC61007FF080C02FFD084402B188C763B184C620319D8C200FFE101805;
defparam spx9_inst_3.INIT_RAM_1E = 288'h3B18401FFC20300BFF421100AC6231D8EC6131880C67630803FF8406017FE84220158C46;
defparam spx9_inst_3.INIT_RAM_1F = 288'h02FFD084402B188C763B184C620319D8C200FFE101805FFA10880563118EC763098C4063;
defparam spx9_inst_3.INIT_RAM_20 = 288'h231D8EC6131880C67630803FF8406017FE84220158C463B1D8C2631018CEC61007FF080C;
defparam spx9_inst_3.INIT_RAM_21 = 288'h319D8C200FFE101805FFA10880563118EC763098C40633B18401FFC20300BFF421100AC6;
defparam spx9_inst_3.INIT_RAM_22 = 288'h06017FE84220158C463B1D8C2631018CEC61007FF080C02FFD084402B188C763B184C620;
defparam spx9_inst_3.INIT_RAM_23 = 288'h63118EC763098C40633B18401FFC20304BFF421100AC6231D8EC6131880C67630803FF84;
defparam spx9_inst_3.INIT_RAM_24 = 288'h1018CEC61007FF080C42FFD084402B188C763B184C620319D8C200FFE101845FFA108805;
defparam spx9_inst_3.INIT_RAM_25 = 288'hC20300BFF421100AC6231D8EC6131880C67630803FF8406417FE84220158C463B1D8C263;
defparam spx9_inst_3.INIT_RAM_26 = 288'h02B188C763B184C620319D8C200FFE101805FFA10880563118EC763098C40633B18401FF;
defparam spx9_inst_3.INIT_RAM_27 = 288'h31880C67630803FF8406017FE84220158C463B1D8C2631018CEC61007FF080C02FFD0844;
defparam spx9_inst_3.INIT_RAM_28 = 288'hFFE101805FFA10880563118EC763098C40633B18401FFC20300BFF421100AC6231D8EC61;
defparam spx9_inst_3.INIT_RAM_29 = 288'h220158C463B1D8C2631018CEC61007FF080C02FFD084402B188C763B184C620319D8C200;
defparam spx9_inst_3.INIT_RAM_2A = 288'h3098C40633B18401FFC20300BFF421100AC6231D8EC6131880C67630803FF8406017FE84;
defparam spx9_inst_3.INIT_RAM_2B = 288'h007FF080C02FFD082402B188C763B184C620319D8C200FFE101805FFA10880563118EC76;
defparam spx9_inst_3.INIT_RAM_2C = 288'h420900AC6231D8EC6131880C67630803FF8406017FE84120158C463B1D8C2631018CEC61;
defparam spx9_inst_3.INIT_RAM_2D = 288'h3B184C620319D8C200FFE101805FFA10480563118EC763098C40633B18401FFC20300BFF;
defparam spx9_inst_3.INIT_RAM_2E = 288'h30803FF8406017FE84120158C463B1D8C2631018CEC61007FF080C02FFD082402B188C76;
defparam spx9_inst_3.INIT_RAM_2F = 288'h0030000CCD63319ACCC663018CCC663019FF420900AC6236341B8C061D8EC6131880C676;
defparam spx9_inst_3.INIT_RAM_30 = 288'h066341B8C061D8EC6131880C676308031A0C66B3318CCC0E33598C666B45B80C66B198CD;
defparam spx9_inst_3.INIT_RAM_31 = 288'hC62331A0DC6031998CC6633188C66633198CC663118763B184C620319D8C200FFB33198C;
defparam spx9_inst_3.INIT_RAM_32 = 288'h061D8EC6131880C67600333198CC66341B8C061D8EC631018CEC61007FD0824C2B331A0D;
defparam spx9_inst_3.INIT_RAM_33 = 288'h420900180C6033FE841260319ACC60B31ACCC68319B8DE6837180CC763018CCC6633198C;
defparam spx9_inst_3.INIT_RAM_34 = 288'hC0233FE04C063198CCC663018763B184C620319D8C200000031BCDD6BB7180CC763019FF;
defparam spx9_inst_3.INIT_RAM_35 = 288'h06E3019FFC2331998C0660318CCC6837180CFFA10498566333190CC063199FF42093FE04;
defparam spx9_inst_3.INIT_RAM_36 = 288'hF619AC43719800EB771018CEC61007FFFE84127FCEC763098C40633B184018D06E30198D;
defparam spx9_inst_3.INIT_RAM_37 = 288'h84422110884422110884422110846231188C46231188C460121108844221108844221108;
defparam spx9_inst_3.INIT_RAM_38 = 288'h84431497C844221108844221108844221108844221108844221108844221108844221108;
defparam spx9_inst_3.INIT_RAM_39 = 288'h600E2793C9E4F2793C9E4F2793C106D211086A420F108846D28908844221108844221108;
defparam spx9_inst_3.INIT_RAM_3A = 288'h9E4F2793C9E4F2793C9E4F2793C9E4F2793C9E4F2793C9E4F2793C6030180C06030180C0;
defparam spx9_inst_3.INIT_RAM_3B = 288'h9E7A2F13C9E4F2793C9E4F2793C9E501B1B09E4F2793C9E4F2793C9E4F2793C9E4F2793C;
defparam spx9_inst_3.INIT_RAM_3C = 288'h16CB4017890590417832594CA0D06894E520B9034003218192ED6506FA2793C844F1593C;
defparam spx9_inst_3.INIT_RAM_3D = 288'h0693CEA0D3BDB01A00069DC1A0A84896E55210480147818192C744B28344B72AB8365B61;
defparam spx9_inst_3.INIT_RAM_3E = 288'hBA56C00653C080F34B96D5A1400848021200310340109365CC1B3184CE260099A4C01330;
defparam spx9_inst_3.INIT_RAM_3F = 288'h324B4006EB79C0B600B41BEE66436CB4BB6E394F0B6643CDCCC86D96976DC729E16EC800;

SPX9 spx9_inst_4 (
    .DO({spx9_inst_4_dout_w[26:0],spx9_inst_4_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[17:9]})
);

defparam spx9_inst_4.READ_MODE = 1'b0;
defparam spx9_inst_4.WRITE_MODE = 2'b01;
defparam spx9_inst_4.BIT_WIDTH = 9;
defparam spx9_inst_4.BLK_SEL = 3'b000;
defparam spx9_inst_4.RESET_MODE = "SYNC";
defparam spx9_inst_4.INIT_RAM_00 = 288'hFF7C411FE000210018007F01000040000000007A0341800000000800868021A880002080;
defparam spx9_inst_4.INIT_RAM_01 = 288'h0000000000000000000000000000000000000000000000010000EE7C000001090080A122;
defparam spx9_inst_4.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_20 = 288'h0B1002C200B0402C08195E0152194CC67341A4D46B361B4EE783C9E8F67C3E9F8FE40062;
defparam spx9_inst_4.INIT_RAM_21 = 288'hB0DA773C1E4F47B3E1F4FC7F200012F80C80054E01D6E091882C480D0183DE60B0002D00;
defparam spx9_inst_4.INIT_RAM_22 = 288'hEB804000CEF1682C001C040017000003F000007A3F440057A0386290CA66339A0D26A359;
defparam spx9_inst_4.INIT_RAM_23 = 288'hECF87D3F1FC800C400FD20015E8F780801E8FD10015E8090010000040039614F6FFBF048;
defparam spx9_inst_4.INIT_RAM_24 = 288'h011E3D7008418803118CC8653319CD069351ACD86D371BCE071391CCE8753B1DCF0793D1;
defparam spx9_inst_4.INIT_RAM_25 = 288'h9CD069351ACD86D371BCE071391CCE8753B1DCF0793D1ECF87D3F1FC80312F800100F1FC;
defparam spx9_inst_4.INIT_RAM_26 = 288'hEB8980418EBED46DD7EC80373C1ECF276BA9406E4C058D0000C4000418A13118CC865331;
defparam spx9_inst_4.INIT_RAM_27 = 288'h2C68000602C00001D9DCF203DD7EB80BAFD94C76731C9D4F64B1D90C7078398E481B9242;
defparam spx9_inst_4.INIT_RAM_28 = 288'h007000818ECEE7CE16ECFE011C00179C01EAECEC7B202EC81001E70C7677214ECEC77260;
defparam spx9_inst_4.INIT_RAM_29 = 288'hECEC772602C68000602C00001C00206373FED8F9FF002E000BCE00F276501FED8F6405D9;
defparam spx9_inst_4.INIT_RAM_2A = 288'hF3863B3B9007000818E8EE7CFF80170005E7000D3A3EA03767B202EC81001E70C7677214;
defparam spx9_inst_4.INIT_RAM_2B = 288'h00773A3B1E880BA200E001031D1DCF9FF002E000BCE001172BB3B1E880BA3D9017640800;
defparam spx9_inst_4.INIT_RAM_2C = 288'hF3F0015E710063C00010060000AE016BBDE7E002BCE0AE000BCFC00579C4018F0000C058;
defparam spx9_inst_4.INIT_RAM_2D = 288'h200C07080EDEFD1680027673BD90576480301C70000200C00015C01079F800AF382B8002;
defparam spx9_inst_4.INIT_RAM_2E = 288'h180E0017B23A0005D9ACF5FB20CEC9006038E000040100C003F40240744002008063C000;
defparam spx9_inst_4.INIT_RAM_2F = 288'h30140B1A000100603840003B34B0BA0009D90FA0011D998F7FBBDBECC8080301C7000040;
defparam spx9_inst_4.INIT_RAM_30 = 288'h00180A0580053E03CD40023B2DFBCF6F81B9DC94373DDE06E77250DCF7F81B9ECEC3B3B9;
defparam spx9_inst_4.INIT_RAM_31 = 288'hD4E050008ECA4E5BDBE06E77250DCF7781B9DC94373DFE06E7B204ECEA763B930140B1A0;
defparam spx9_inst_4.INIT_RAM_32 = 288'hDCEE4A1B9EEF0373B9286E7BFC0DCF640DD9D4EC7726028163400030140B0007EABFE7B1;
defparam spx9_inst_4.INIT_RAM_33 = 288'h9000080301C0023DE84077FBE80200C071C000180A0580017F47B1D4CC50008EC90FB7C0;
defparam spx9_inst_4.INIT_RAM_34 = 288'h94D8035E1EC8BA00046C7265228ECF267206E196B92989C83A721290C8653319CB81A0D8;
defparam spx9_inst_4.INIT_RAM_35 = 288'h0970782800258031E1FF7441DD9E88EBA298CD76A31D9ECCC7B1C9EC80BB3C98001135C9;
defparam spx9_inst_4.INIT_RAM_36 = 288'h03053BE18DC980A058D0001C0D06C20101C6E8F47FDD1A5A0380AEE070415C030703820C;
defparam spx9_inst_4.INIT_RAM_37 = 288'h208E46229108642209CCA00E078A0000C0502C20101E2EFF7C01B9DC80B73194077E3E1A;
defparam spx9_inst_4.INIT_RAM_38 = 288'h0074400000C0C00044AB29B6C000C66405D9E480AE44AE3F1C0018CCF6731D9E8EE773C8;
defparam spx9_inst_4.INIT_RAM_39 = 288'hECF4411D144A03921440003A334EC80BB3D1047450E80E0003A34CEC80BB3D104746DA80;
defparam spx9_inst_4.INIT_RAM_3A = 288'hE8B83B202ECF4411D128A03921040003A2FCEC80BB3D104744DA80E48500400E8C63B202;
defparam spx9_inst_4.INIT_RAM_3B = 288'hEC80BB3E9252A3B202ECF4411D10CA03922040003A2C4EC80BB3D1047446A80E48110000;
defparam spx9_inst_4.INIT_RAM_3C = 288'h000633202ECBB0C0000C66405D9EC80BB3C90C6800018CC80BB2180A7243DC9EC80BB29C;
defparam spx9_inst_4.INIT_RAM_3D = 288'h390003199017655C60000633202ECF6405D9E486340000C66405D90C053921EE4B779472;
defparam spx9_inst_4.INIT_RAM_3E = 288'hDC980B1A000300E07840200C4000C667B3D9017668E80E3D3434060A71C2400AD9293FCA;
defparam spx9_inst_4.INIT_RAM_3F = 288'h066E405B9036E780FEE001B7202DC80015B9026537206DCF013100E001B7206036E7A3DF;

SPX9 spx9_inst_5 (
    .DO({spx9_inst_5_dout_w[26:0],spx9_inst_5_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[17:9]})
);

defparam spx9_inst_5.READ_MODE = 1'b0;
defparam spx9_inst_5.WRITE_MODE = 2'b01;
defparam spx9_inst_5.BIT_WIDTH = 9;
defparam spx9_inst_5.BLK_SEL = 3'b001;
defparam spx9_inst_5.RESET_MODE = "SYNC";
defparam spx9_inst_5.INIT_RAM_00 = 288'h000204018F0000803800003AFD9FC103800AEC803AE80EC90071C000180B000EF8037204;
defparam spx9_inst_5.INIT_RAM_01 = 288'h1C70000200C001100210063C00010060008210063C0001006000000408031E0000803000;
defparam spx9_inst_5.INIT_RAM_02 = 288'hE8863D7D10C764B1FE0780021EBE8F64A1B91A6E772602C68000401C001040641767B240;
defparam spx9_inst_5.INIT_RAM_03 = 288'h0077C5C00047A37E803016340003016000002D3F811EB00023D6120040011EB00023D600;
defparam spx9_inst_5.INIT_RAM_04 = 288'hEF80373B9016E77280EFEFC34060A77C31B930140B1A000180B000006FFD1F8020105DDF;
defparam spx9_inst_5.INIT_RAM_05 = 288'hE4CA451D9E4CE40D7B2D7253139074E4252190CA6633970341B12000180A05840203C5DF;
defparam spx9_inst_5.INIT_RAM_06 = 288'hE883BB3D11D745319AED463B3D998F6393D90176793000226B9329B006BC3D91740008D8;
defparam spx9_inst_5.INIT_RAM_07 = 288'h00381A0D8402038DD1E8FFBA303407015DC0E082B8060E07041812E0F050004B0063C3FE;
defparam spx9_inst_5.INIT_RAM_08 = 288'hCC80BB3C9015C895BFDF8003199ECF03B3D1D8EC790411C8C452210C8441399401C0F140;
defparam spx9_inst_5.INIT_RAM_09 = 288'h01767A208E89DD01C00074699D901767A208E8AF50000E88000018340008956536D80018;
defparam spx9_inst_5.INIT_RAM_0A = 288'h00745F9D901767A208E8A9501C90A00801D18C76405D9E8823A2C14072428800074669D9;
defparam spx9_inst_5.INIT_RAM_0B = 288'h4072440800074589D901767A208E89B501C90220001D17076405D9E8823A289407242080;
defparam spx9_inst_5.INIT_RAM_0C = 288'h017679218D00003199017643014E487B93D90176539D901767B24A5476405D9E8823A251;
defparam spx9_inst_5.INIT_RAM_0D = 288'hEC80BB3C90C6800018CC80BB2180A7243DC96EF28E4000C66405D9761800018CC80BB3D9;
defparam spx9_inst_5.INIT_RAM_0E = 288'h2D07BB226ECCDD01BF9E8680C14DF848014B2527F9472000633202ECAB8C0000C66405D9;
defparam spx9_inst_5.INIT_RAM_0F = 288'h200E38000601C0F080400E80018CCF67B202ECFCB83FEE080000000002B82660006A0004;
defparam spx9_inst_5.INIT_RAM_10 = 288'hECF6480301C70000200C002BC2010063C00010060015E1008031E0001007080ECF6461D9;
defparam spx9_inst_5.INIT_RAM_11 = 288'h0A26001B9046E41C00DC8237208DCA0333B930140B1A000100603800003B280DA823B200;
defparam spx9_inst_5.INIT_RAM_12 = 288'hECF673E80E482B0680E4D97A3C9ECEE4C0502C6800060281610018046E531D9006E7B3FE;
defparam spx9_inst_5.INIT_RAM_13 = 288'h400610000ECF6480301C7000040180E001BD4011BB3D9200C071C000180A0580057FE9B9;
defparam spx9_inst_5.INIT_RAM_14 = 288'h03003B202EC843A3D9200E38000200C07000E7A0031D0ECF6480301C7000040180E0019D;
defparam spx9_inst_5.INIT_RAM_15 = 288'hEC80031EBE8F6772602C68000401C2013000E8F47FDD140003B3E60074405D1007644480;
defparam spx9_inst_5.INIT_RAM_16 = 288'hE881373C01F700C1D1036E7803EE076411B9E007B804AEC82B73C07F700A5D9E880021EB;
defparam spx9_inst_5.INIT_RAM_17 = 288'hEC82005D904023B2080C023B3D9200E38000301600000DCF00FDC02474405B9E01FB8054;
defparam spx9_inst_5.INIT_RAM_18 = 288'h3C003B2982A70200046C1E005D93070200046C0C009D900003D606017641006EC8207C06;
defparam spx9_inst_5.INIT_RAM_19 = 288'h1F01BB2982570200046C06811D92902BB200087AD35C080011B4C8067653048E040008D8;
defparam spx9_inst_5.INIT_RAM_1A = 288'hD000080301C00263D103307A208EFF7FA280200C071C00010070000000011EB00063D698;
defparam spx9_inst_5.INIT_RAM_1B = 288'h1A20139EB40663B202407AC90802E7AD0018CC7640480F586363D9DC8D07DB9D8EE4C058;
defparam spx9_inst_5.INIT_RAM_1C = 288'h3016340003016000A04E7AD0198EC80941EB0A280B9EB4006331D901283D618D8F6781B9;
defparam spx9_inst_5.INIT_RAM_1D = 288'hE06E468884E7AD0198EC80911EB24220B9EB4006331D901223D618D8F6772341F6E763B9;
defparam spx9_inst_5.INIT_RAM_1E = 288'h007A84018F0000C058002A139EB40663B202547AC28A82E7AD0018CC76404A8F586363D9;
defparam spx9_inst_5.INIT_RAM_1F = 288'h047AC0008F5800B5FEFF823D600047AD4018D8F6763B9301634000100600000E0023D5C0;
defparam spx9_inst_5.INIT_RAM_20 = 288'hD88237200DCA6001B1006E421B94C0036210DC84021B92C06001B1086E42808D88013400;
defparam spx9_inst_5.INIT_RAM_21 = 288'h0C6E53000D88637208DC9603000D88237212046E53000D88237212010436208DC9603000;
defparam spx9_inst_5.INIT_RAM_22 = 288'hE0000803800063B210017641002EC803B3D9200E38000301600000DC9603000D88037212;
defparam spx9_inst_5.INIT_RAM_23 = 288'h200E000604D767D6600C764D154AD7AFB2401C70000401C00031D94C74431D9E8F648038;
defparam spx9_inst_5.INIT_RAM_24 = 288'hECC00089AE88036204206E7A2003D76763B930140B1A000080300034552B5EB10063C000;
defparam spx9_inst_5.INIT_RAM_25 = 288'hDC82019B1026E7809880701300ED8F01300CD88236202DCF00A1D9006E781D9ECFF889D9;
defparam spx9_inst_5.INIT_RAM_26 = 288'h077641804EC828A9D904103B200A0007B3D9200E3800030140B0008F7A41DB9056C41008;
defparam spx9_inst_5.INIT_RAM_27 = 288'hE0000803800023B3C02C5FB8008EC84811D9E02038008EC84BA3D1EC90071C0001007000;
defparam spx9_inst_5.INIT_RAM_28 = 288'hE072781D14D76793D1EC9006038E000080301C0001020F481BAFD961767AE80EC9006038;
defparam spx9_inst_5.INIT_RAM_29 = 288'h2400101D7EB80BAE14EA993B3D54075D0080EC9006038E000080301C00011D9E01038098;
defparam spx9_inst_5.INIT_RAM_2A = 288'h046E411DF046E772602C6800040180E00008907A40DD7ECD4C60004075FAE58FE75C2967;
defparam spx9_inst_5.INIT_RAM_2B = 288'h281634000301600008DCF0011C0046E42008EFF7C11B9DC980B1A000180B000FB013BFDF;
defparam spx9_inst_5.INIT_RAM_2C = 288'hE0023D375F4C8FD2804077D7A080020101BBEFF7E81C0E013B7BBDFF6F77680DEA010060;
defparam spx9_inst_5.INIT_RAM_2D = 288'h40FA501BB38CA000081770011E9A3FA53BE9407037A8FE400101BDDEFFB7A9FF0000102E;
defparam spx9_inst_5.INIT_RAM_2E = 288'hE013B7BBDFF6F77A8030140B1A000180A05800447D231F4808AAB8000205DC0047A657E9;
defparam spx9_inst_5.INIT_RAM_2F = 288'hDEEF7FDBDF8EE00080DEFEF9000040BB8008F4B47D27FF4A0101DF0C8200080EFF7E81C0;
defparam spx9_inst_5.INIT_RAM_30 = 288'hF484101AF4C000102EE0023D285F48CFD2800177F9B10000205DC0047A547E9FCFA501C0;
defparam spx9_inst_5.INIT_RAM_31 = 288'h007D005D9EC80021EC057640010F60000010F610071C000180A05840777BA06F49A7D3E7;
defparam spx9_inst_5.INIT_RAM_32 = 288'hD48036208F6000B5FEFFEE7D9F401767B200087B015D900043D9A9D8EE4C058D00008038;
defparam spx9_inst_5.INIT_RAM_33 = 288'h2C7F8005E02765306001764E000ECF648038E0000C058000000410F60280006087B01802;
defparam spx9_inst_5.INIT_RAM_34 = 288'h4C161806C01764E000ECF648038E000080380000021EB4C07811D94C16000002801BB298;
defparam spx9_inst_5.INIT_RAM_35 = 288'h0017809D930003B3D9200E38000200E000000C7AD3408ECA6000500376530581F98009D9;
defparam spx9_inst_5.INIT_RAM_36 = 288'h01043B298021081DD94C7F8900CECA6000500576530002B023B2982C000B006ECA60B1FE;
defparam spx9_inst_5.INIT_RAM_37 = 288'h200E000002D7F811EB00023D6120000011EB00023D612ECF648038E0000803800003D698;
defparam spx9_inst_5.INIT_RAM_38 = 288'h0006201EB40113BBDD4010071C0001007080E07FB80000C203D68022777BA80200E38000;
defparam spx9_inst_5.INIT_RAM_39 = 288'hE000040180000005EB007AC4018F000040180000009EB007AC4018F0000803840703FDC0;
defparam spx9_inst_5.INIT_RAM_3A = 288'h1C70000401C000009C0D203D6802277D0070EEFF80018407AD0044EFF7501DF402008038;
defparam spx9_inst_5.INIT_RAM_3B = 288'h281634000200E000004C06901EB40113BFFE0006201EB40113BE8038777BA80EFA010040;
defparam spx9_inst_5.INIT_RAM_3C = 288'hE9883A2A0CFA0100703C60000602816001EA0B777BA02EEEA50080DFF03BA14EEEFD0060;
defparam spx9_inst_5.INIT_RAM_3D = 288'hDA81B6606D8EBC0DAD016A7FDBF4070793FEE38438A10E1F040D8F40747B202EB80BAA02;
defparam spx9_inst_5.INIT_RAM_3E = 288'h401B501C0EC87BB2A048262C000401C0F0001880AC280CFFE80400F5801BBE3406A773B7;
defparam spx9_inst_5.INIT_RAM_3F = 288'hF205BB3D901767EAA8002032018F0913B21AEC82E9000F005BB3D9017672018F0913B280;

SPX9 spx9_inst_6 (
    .DO({spx9_inst_6_dout_w[26:0],spx9_inst_6_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[17:9]})
);

defparam spx9_inst_6.READ_MODE = 1'b0;
defparam spx9_inst_6.WRITE_MODE = 2'b01;
defparam spx9_inst_6.BIT_WIDTH = 9;
defparam spx9_inst_6.BLK_SEL = 3'b010;
defparam spx9_inst_6.RESET_MODE = "SYNC";
defparam spx9_inst_6.INIT_RAM_00 = 288'h0C7B40008EC843DA00047B401EDEC90071C00028120980074CF0004075FAE1EE000011EB;
defparam spx9_inst_6.INIT_RAM_01 = 288'hF68C3B200F680135ED1076401ED0070005EAE0003D41014764009AF68A3B200F680021D9;
defparam spx9_inst_6.INIT_RAM_02 = 288'hEC8420001EC820FC00EC88011D914013B2300176400003D767B2401C70000401C000009A;
defparam spx9_inst_6.INIT_RAM_03 = 288'h0E767B2401C70000401C00001FCF6803DA0C0000BDA00F683BB3D9200E38000200E00018;
defparam spx9_inst_6.INIT_RAM_04 = 288'h2C68000401C00001C02D7F3D5C0007A801FAF6803DA1C0070005EAE0003D400027B401ED;
defparam spx9_inst_6.INIT_RAM_05 = 288'hF57000006F500135D9F6803DBD9200E380003016101D9EC813B202041637200F6F677260;
defparam spx9_inst_6.INIT_RAM_06 = 288'hEC90071C000100603800032D1FF4077C0002C87FFBE80200C071C0001007000007000406;
defparam spx9_inst_6.INIT_RAM_07 = 288'hEC88811D91076441D901083B218EC81811D90C76431D901063B200EB86831D900767AE80;
defparam spx9_inst_6.INIT_RAM_08 = 288'h281634000200E10000E8F648038E0000803800043B2060476421D9087640410EC883B208;
defparam spx9_inst_6.INIT_RAM_09 = 288'h0076405D9B8DE00080400003048ECF600002EC88BB38FE8001AC48026E41402DCEC77260;
defparam spx9_inst_6.INIT_RAM_0A = 288'h2476500001A200F3D1400003048ECB600050ECF4411B14E729009B8800100000C123B368;
defparam spx9_inst_6.INIT_RAM_0B = 288'h002000018247674000EC80BB22080F4000804020030182476440000806091D9280000018;
defparam spx9_inst_6.INIT_RAM_0C = 288'hC0000C0502C2010000022EE20000530DE0000920022E8002000018247668000CE2005348;
defparam spx9_inst_6.INIT_RAM_0D = 288'hE880000000002BA266002549000F9767FDD9000000000057671C1C0002811E881A00E078;
defparam spx9_inst_6.INIT_RAM_0E = 288'hE09980049A400011994110FE5C9FF72400000000015C933000DFC80068743D8007CBA3FE;
defparam spx9_inst_6.INIT_RAM_0F = 288'h0130C0402F96E7FDB9000000000056E4CC0011B200080C8E4421F2E0FFB820000000000A;
defparam spx9_inst_6.INIT_RAM_10 = 288'h01203E5A9FF6A400000000015A9E403A3202017CB63FED880000000002B63C8076CD7A28;
defparam spx9_inst_6.INIT_RAM_11 = 288'hBF2000008D898005774C0001806DC82005B9D8EE4C0502C68000200C20100200C7838AFB;
defparam spx9_inst_6.INIT_RAM_12 = 288'h407000018E4F666BD00020031C9EC8401DD917767A280B32000010D8843A2020401373C9;
defparam spx9_inst_6.INIT_RAM_13 = 288'h33009DAD8000300DB90400B73B1DC980A058D0000C0502C20101D0E8F67B202ECC8F4000;
defparam spx9_inst_6.INIT_RAM_14 = 288'hFC0010018E4A0089D90A01BB234ECF4500DC4000021B1087440408026E792F44000011B1;
defparam spx9_inst_6.INIT_RAM_15 = 288'h0601B73B1DC980A058D0000C0502C20101CAE8F67B202ECA4F80004000031C940113B2A7;
defparam spx9_inst_6.INIT_RAM_16 = 288'hDC980A058D0000C0502C2010000EBF67AE802F2000010D8F64D4800002362240118E2000;
defparam spx9_inst_6.INIT_RAM_17 = 288'h2C680006028161008000747B3D10B2000010D8F6444800002362220106C60000601B73B1;
defparam spx9_inst_6.INIT_RAM_18 = 288'h5974421C901030C000DC86BA220E481018B00000B720C7800005B91018001B9ECEE4C050;
defparam spx9_inst_6.INIT_RAM_19 = 288'hECE8031C10C747B21239704305EE0A18C410E882841D137053A3C10006393B95574429C9;
defparam spx9_inst_6.INIT_RAM_1A = 288'h94AA0000AECE4831C10C747B212467043080E089BB3520C70431D1EC84999C10C3038242;
defparam spx9_inst_6.INIT_RAM_1B = 288'h2C203B3500006393B9E480B9200808E00008ECE8031C10C747B212E0983A21A2F704502A;
defparam spx9_inst_6.INIT_RAM_1C = 288'h980023FD163A000010D8F65A6800002362320132F10000601B73B1DC980A058D0000C050;
defparam spx9_inst_6.INIT_RAM_1D = 288'h002000010F59CDC00040003D67F7C00080301C70000602816100804CCC0013FECF4404A7;
defparam spx9_inst_6.INIT_RAM_1E = 288'h0076500800006201EB40113B2000C203D6802276461D928B4000576000100000C7ACCAD0;
defparam spx9_inst_6.INIT_RAM_1F = 288'h402001280E076435D9FC9C001FFFC00080301C7000040180E10080E705BB3D9017644A60;
defparam spx9_inst_6.INIT_RAM_20 = 288'h1C20101E40B767B202ECEEF1000402000E80E076435D9E8FC001E40B767B202ECF8C5000;
defparam spx9_inst_6.INIT_RAM_21 = 288'h00043636F5C0024802BCAC0000C036E45C8066B8000800002363B1DC980A058D00008030;
defparam spx9_inst_6.INIT_RAM_22 = 288'hD8B61E3AF98FC0000EE01638002026E780024023C90004000011B18328501DDEEA02F680;
defparam spx9_inst_6.INIT_RAM_23 = 288'hEFF7C05DFC4A0101DFED84BBE1E036E7B6808FA000010D8C4F500031200C3C0002000008;
defparam spx9_inst_6.INIT_RAM_24 = 288'h407BCE0004000011B1340097A70001C2BA804077FB7DF403A500000C6C43808DCA43D816;
defparam spx9_inst_6.INIT_RAM_25 = 288'hEF8238058E000809B9E000901C3F80010000046C474F748860000CE01638002026E78002;
defparam spx9_inst_6.INIT_RAM_26 = 288'h9BA0222800A01AF2370C002E37950241316000180A0584020008022CE20005FC0000245D;
defparam spx9_inst_6.INIT_RAM_27 = 288'h3F003A3B1227653680C8F24268000062E3D10FA000010B8F64568000022E24E0108C0000;
defparam spx9_inst_6.INIT_RAM_28 = 288'h54000420E016E76AA0006E763B930140B1A0002812098402001E80C8E8430003D7273218;
defparam spx9_inst_6.INIT_RAM_29 = 288'hEC0001804DCEC7726028163400030140B080400850018F828BB3D9D7A000008D887005A7;
defparam spx9_inst_6.INIT_RAM_2A = 288'h0074467D108013B2309CDE001D115F442002ECF46C6800004363D9B7A000008D89780567;
defparam spx9_inst_6.INIT_RAM_2B = 288'h749A001B9D8EE4C0502C680006028161008084980000888BE001D11FF442006EC8724B38;
defparam spx9_inst_6.INIT_RAM_2C = 288'hEFA0080301C7000060281610080E6DC7B3D96FA000008D885804D73400316800800B7337;
defparam spx9_inst_6.INIT_RAM_2D = 288'h04003300038CE000B15CD829150AC2800040180E1001EEF81BFC97CC0001872EF820BDDF;
defparam spx9_inst_6.INIT_RAM_2E = 288'h000216330400CE50001CBC0003F580008A9000079019340201E200042C613017CBC43010;
defparam spx9_inst_6.INIT_RAM_2F = 288'h9BA000002EC8602880A3A0001D9E886163D9082C61C0208C60000C042E6A080B2A0100F9;
defparam spx9_inst_6.INIT_RAM_30 = 288'h7BA00000EEC860288083A00000CECF0432808BA000008EC860288093A000006ECF243280;
defparam spx9_inst_6.INIT_RAM_31 = 288'h402E50000047443014403250000037476219403650000017443014403A50000E8EE43280;
defparam spx9_inst_6.INIT_RAM_32 = 288'hDC82009C1106E4483EDC8AB822E0C7074219402650000077443014402A50000067475219;
defparam spx9_inst_6.INIT_RAM_33 = 288'hDCB9781B171F0352E1E0687FC0280C00000CCCE65000401018F1A1041E3520E186C4283A;
defparam spx9_inst_6.INIT_RAM_34 = 288'h082C75C0258E60000C042E6488002A0101010002163D0C1A0100E175F0392E9E0705CFC0;
defparam spx9_inst_6.INIT_RAM_35 = 288'hDBA000008C88602880E3A000006C8E043280EBA000002C88602880F3A000191C48616391;
defparam spx9_inst_6.INIT_RAM_36 = 288'h405E5000004624301440625000003626E219406650000016243014406A50000C4DE43280;
defparam spx9_inst_6.INIT_RAM_37 = 288'hBC8200981105E4483EBC8AB022E0C606C219405650000076243014405A5000006626D219;
defparam spx9_inst_6.INIT_RAM_38 = 288'hBCB57817169F02D2D1E05857C02E0800000CACD65000401018F161041E2D20E185C4283A;
defparam spx9_inst_6.INIT_RAM_39 = 288'h015614400A8F02B06000546A3954000020B122201A28040424000858A7100D9E0605AFC0;
defparam spx9_inst_6.INIT_RAM_3A = 288'h63CC5933965F94048060CEC9000040097248405043D51A4922A2580156D10000670131C0;
defparam spx9_inst_6.INIT_RAM_3B = 288'hD8EE4C0502C6800160A4542B0804040F700090C66230FE0002733194C45831961C858B29;
defparam spx9_inst_6.INIT_RAM_3C = 288'hDC980A058D0000C0502C20101B5ECF65B6800002362140134F3000FA83805B970E4001B9;
defparam spx9_inst_6.INIT_RAM_3D = 288'hD89AE400031008EA480003011B9D8EE4C0502C6800060281610000E5FA501D12AA03A3B1;
defparam spx9_inst_6.INIT_RAM_3E = 288'hB400101DBEA8B1302CEE8B09DDFEDA00B6800006363DD401A50000086C7BE803BA000008;
defparam spx9_inst_6.INIT_RAM_3F = 288'hD893005EF5C0001806DCEC7726028163400030140B0804049D0080EAF6C3B5800203AA27;

SPX9 spx9_inst_7 (
    .DO({spx9_inst_7_dout_w[26:0],spx9_inst_7_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[17:9]})
);

defparam spx9_inst_7.READ_MODE = 1'b0;
defparam spx9_inst_7.WRITE_MODE = 2'b01;
defparam spx9_inst_7.BIT_WIDTH = 9;
defparam spx9_inst_7.BLK_SEL = 3'b011;
defparam spx9_inst_7.RESET_MODE = "SYNC";
defparam spx9_inst_7.INIT_RAM_00 = 288'h4072F9680B9A039BCD4C703FDC0E8F00B100007009DC0ECF47D6800004363D9FBA000008;
defparam spx9_inst_7.INIT_RAM_01 = 288'h02744280EECF4716800004323D9CBA000008C8E473280381E3000030140B0804068FA000;
defparam spx9_inst_7.INIT_RAM_02 = 288'hF5978052F8C0026A78004ECB0000C7277280AFA000018C8F25000401018119904013320E;
defparam spx9_inst_7.INIT_RAM_03 = 288'hFF6E5DA3800200B018167078200707AC00006C7AC00D8F580035D96C7AC91D11E0000008;
defparam spx9_inst_7.INIT_RAM_04 = 288'h4A0095B580003009B9D8EE4C0502C6800080381E100800016BFDFF047AC0008F5F1373B9;
defparam spx9_inst_7.INIT_RAM_05 = 288'h2D7F9FFEB007ACAC300276415D90F00BB25E02764009A017AC01EB07767B2B54000011B1;
defparam spx9_inst_7.INIT_RAM_06 = 288'h0003000004D403D600F5800B5FE7FFAC01EB150013400F5803D6002D7F9FFEB007AC8C00;
defparam spx9_inst_7.INIT_RAM_07 = 288'hECC0000201879801FE0879801FE0479880301C70000602816100800000011EB060084B98;
defparam spx9_inst_7.INIT_RAM_08 = 288'hE8BFBB3D1047440000E8A003100E885BA3D900003CDCF34001E2004D003CC58FF00FB258;
defparam spx9_inst_7.INIT_RAM_09 = 288'hE8DADC000040003100E8803A21CE8F6461D98069A05D9ECC03B2004D003CC58FF00FB3E6;
defparam spx9_inst_7.INIT_RAM_0A = 288'h1900A5A000003009B9D8EE4C0502C6800040180E10080E740BB3D980767C1D17F767A208;
defparam spx9_inst_7.INIT_RAM_0B = 288'h28163400030140B0804001004FFA400018D9F402009D90C397D00801767B3354000011B1;
defparam spx9_inst_7.INIT_RAM_0C = 288'h060133391CCA00E078C0000C0502C20000C74C00101DDEEA0166082079C00A4F3EC77260;
defparam spx9_inst_7.INIT_RAM_0D = 288'hECEC5001880063B3C1107678250E892BA3B90022FF000E0F2556800002322740128C4000;
defparam spx9_inst_7.INIT_RAM_0E = 288'h3C201002F5800369B9E8F4405D14DA0362000C707924F94003BDFEECF6405D9007000018;
defparam spx9_inst_7.INIT_RAM_0F = 288'hE89ABA3B9007CFF000E0F2426800002322940102C5000060133391CCA00E078C00010070;
defparam spx9_inst_7.INIT_RAM_10 = 288'h80063B3C14000031D9D888B80000C40031D9E080031D9D8903B283406C40018E0F278250;
defparam spx9_inst_7.INIT_RAM_11 = 288'hD000100703C2010177E800329B9E8F4405D1C484001BEFF767B202EC83B3AC0002010018;
defparam spx9_inst_7.INIT_RAM_12 = 288'h2C20101414006003D9A5F667BB800766B6800002362240154FB0000601373B1DC980A058;
defparam spx9_inst_7.INIT_RAM_13 = 288'h7DA003001E4C1792F7AC00101BDDEA01C6082079C00A4F3F079391CCA00E078C0000C050;
defparam spx9_inst_7.INIT_RAM_14 = 288'hE0F27BDFEECF6405D9007000018ECEA5001880063B3C1107678250E892BA3B10038CE000;
defparam spx9_inst_7.INIT_RAM_15 = 288'hD480031C1E4F04A1D135747620040CA000879000369B1E8F4405D14C94000F9406A40018;
defparam spx9_inst_7.INIT_RAM_16 = 288'h070ADF0004020031000C767828000063B3A911700001880063B3C100063B3A9207662280;
defparam spx9_inst_7.INIT_RAM_17 = 288'h107AC0880200C071C000200E078402000B600065363D1E880BA217240037DFEECF6405D9;
defparam spx9_inst_7.INIT_RAM_18 = 288'h180E38000200C070800069C81EB40707B202E880B9202E0810108B407071A30F58410197;
defparam spx9_inst_7.INIT_RAM_19 = 288'h08766DB20006C77260281634000301610080ECEC772602C6800040180E10080D5F47B240;
defparam spx9_inst_7.INIT_RAM_1A = 288'h007646DD9F1003B3D90476400004006001D94006003D90E767DC00ECF6411D90006001D9;
defparam spx9_inst_7.INIT_RAM_1B = 288'h2C20100000072001D9EC823B2FFC8003B280400003001EC8003000EC878001800F640018;
defparam spx9_inst_7.INIT_RAM_1C = 288'h549A000302C00040100C780002008060019F207AC04CF800004CC0000802018F0000C050;
defparam spx9_inst_7.INIT_RAM_1D = 288'h1004031E00008020180054C81EB0420FA0001D7C0002008063C000100403000BC903D604;
defparam spx9_inst_7.INIT_RAM_1E = 288'h080600107207AC4037500009D20000802018F000040100C0025A40F5840BB38001131000;
defparam spx9_inst_7.INIT_RAM_1F = 288'h407AEE00031140002008063C00010040300070903D6400882000585C00040100C7800020;
defparam spx9_inst_7.INIT_RAM_20 = 288'h000802018F000040100C0012A40F5C038AD8001BBD0001004031E0000802018002EC81EB;
defparam spx9_inst_7.INIT_RAM_21 = 288'h10040300024903D600BCEA000848C00040100C780002008060006F207AC019F20000F180;
defparam spx9_inst_7.INIT_RAM_22 = 288'hF58025A780027090001004031E00008020180008C81EB0054E2000482C0002008063C000;
defparam spx9_inst_7.INIT_RAM_23 = 288'hBC00040100C78000200806001D7207AC0107F00014DE0000802018F000040100C003FA40;
defparam spx9_inst_7.INIT_RAM_24 = 288'h0008020180062C81EB002ED60005E440002008063C000100403000D8903D60070D2000B0;
defparam spx9_inst_7.INIT_RAM_25 = 288'h207AC026FC0001AC40000802018F000040100C002CA40F58012A180032150001004031E0;
defparam spx9_inst_7.INIT_RAM_26 = 288'h775C0002008063C0001004030008C903D60224BA000E2EC00040100C780002008060013F;
defparam spx9_inst_7.INIT_RAM_27 = 288'hF000040100C0019A40F5823FBB8003EA10001004031E0000802018003CC81EB0208CA000;
defparam spx9_inst_7.INIT_RAM_28 = 288'h40903D620D8A2001101C00040100C78000200806000A7207AC21D7900020CA0000802018;
defparam spx9_inst_7.INIT_RAM_29 = 288'h0049AD0001004031E00008020180016C81EB2062FE0008D740002008063C000100403000;
defparam spx9_inst_7.INIT_RAM_2A = 288'h0C780002008060000F207AE013F600026500000802018F000040100C0006A40F5A02CB58;
defparam spx9_inst_7.INIT_RAM_2B = 288'h0070C81EB003CF2000A50C0002008063C000100403000F4903D6008C8A0013E4C0004010;
defparam spx9_inst_7.INIT_RAM_2C = 288'h30002C560000802018F000040100C0033A40F58019AF80055B90001004031E0000802018;
defparam spx9_inst_7.INIT_RAM_2D = 288'h08063C000100403000A8903D60040F2001707C00040100C7800020080600177207AC00A7;
defparam spx9_inst_7.INIT_RAM_2E = 288'h0C0020A40F58006A980062050001004031E0000802018004AC81EB0016E6000BE2400020;
defparam spx9_inst_7.INIT_RAM_2F = 288'h1076401D12C727A3C900103D7D10C103D607F0003C1A0000020078F59006038E00004010;
defparam spx9_inst_7.INIT_RAM_30 = 288'hF58000278F59006038E000080301C003BC3EECF6405D9000003044ECD20001001763B3D1;
defparam spx9_inst_7.INIT_RAM_31 = 288'h047AC00023C7AFB61EE000011EBEEFFB806000023D640180E38000200C070005EF640008;
defparam spx9_inst_7.INIT_RAM_32 = 288'hF59006038E000080380077C0004F40000878F590071C00010060380056F800040774001E;
defparam spx9_inst_7.INIT_RAM_33 = 288'h400003C00047ADEA680000000187000089D91C083B2002D3E0F1EB00023D7D91F1980008;
defparam spx9_inst_7.INIT_RAM_34 = 288'h0620006000A00BBFDF0002BD440180E38000200C0700000010005AFF7FC11EB00023D6E7;
defparam spx9_inst_7.INIT_RAM_35 = 288'h0801BD4194076FB600F405821DF000200DEA44E800080EEF7401E80D023BE9FD40004200;
defparam spx9_inst_7.INIT_RAM_36 = 288'h07000629C4D26171B0000802018002DC8AB80033C40100C7800040180E00000FF01BD400;
defparam spx9_inst_7.INIT_RAM_37 = 288'h0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F;
defparam spx9_inst_7.INIT_RAM_38 = 288'h078381C0E0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F;
defparam spx9_inst_7.INIT_RAM_39 = 288'h0984C26130984C26130984C2613098381E0F0703C1C0F078381C0F0783C1E0F0783C1E0F;
defparam spx9_inst_7.INIT_RAM_3A = 288'h0984C26130984C26130984C26130984C26130984C26130984C26130984C26130984C2613;
defparam spx9_inst_7.INIT_RAM_3B = 288'h0984824130984C26130984C26130984824120984C26130984C26130984C26130984C2613;
defparam spx9_inst_7.INIT_RAM_3C = 288'hDBA5801120F0C02D125CABD760502C6020309801400BC5E4C864B10284826130904C2413;
defparam spx9_inst_7.INIT_RAM_3D = 288'h428AC6F851B8D10A00428DC0A00090F03C3002EC220105E4CB653218014781E180152DB1;
defparam spx9_inst_7.INIT_RAM_3E = 288'h170C800BC0006170B24B0C24200C9002240055E140012004CA0A180C0113718022663004;
defparam spx9_inst_7.INIT_RAM_3F = 288'h0865801325B0416800190E473321C05800BA0F8C0641A5D0E664380B001741F182C83000;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[29:0],sp_inst_8_dout[19:18]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[19:18]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b01;
defparam sp_inst_8.BIT_WIDTH = 2;
defparam sp_inst_8.BLK_SEL = 3'b000;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000021C06DF304B000300000A1;
defparam sp_inst_8.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_08 = 256'hFFC0C3C3C3040CFDC050028C3C38FFFFFFFFFC2021222100000033FFFFFFFFF0;
defparam sp_inst_8.INIT_RAM_09 = 256'h3003F3CF77F77DCCC2F3CFFF70C00FFFFFFFFFFFFFFFCDA30CC3FFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_0A = 256'h3FCC43FC4C3FCF30CF10FF130F3CC33CFC30010FFC4CF7F310FCF133FCC33CFC;
defparam sp_inst_8.INIT_RAM_0B = 256'h03004FD3D3FFF03003D3FCC0C00C700C01FD3F30300134C4D30C005F4C4D30C0;
defparam sp_inst_8.INIT_RAM_0C = 256'hC0077D03003BE4FDF7DF7DF3FC0C00FBE4FF7DF7DF7CFF03003E4FF7DF7DF7FF;
defparam sp_inst_8.INIT_RAM_0D = 256'h0000C0C017F3CF7C0CC0C017FFD4711C3D33F3CD03FFCF83F3C83CFCCCCCFFC0;
defparam sp_inst_8.INIT_RAM_0E = 256'hCE0CF3DC4CCF3DC4CCF3DC4CCF3DC0CCF3DC4CCF3D4CCF3D30300C33C0F0F3FF;
defparam sp_inst_8.INIT_RAM_0F = 256'h33344CC33CD74C3FC3005C3F39E0308F033C0CF3CC33CCFC0CF033CF30CF33CC;
defparam sp_inst_8.INIT_RAM_10 = 256'h303D0C00630C130CCF3703F33C30003C30000C000C00030000C00FC4CDC300CC;
defparam sp_inst_8.INIT_RAM_11 = 256'h005FFF51C470F4CFCF340FFF3E0FCF20F3F33333FF03005FCF3DF03303003F03;
defparam sp_inst_8.INIT_RAM_12 = 256'h71333CF71333CF71333CF70333CF71333CF5333CF4C00030CF03C3CFFC000303;
defparam sp_inst_8.INIT_RAM_13 = 256'h0C0170FCFFC00F080CE780C23C0CF033CF30CF33F033C0CF3CC33CCF333833CF;
defparam sp_inst_8.INIT_RAM_14 = 256'h7CF030034F03003FFDCDFFF03004333F0330CCDF03000DCCF030000C000301F3;
defparam sp_inst_8.INIT_RAM_15 = 256'hC30C0F0C00D17345CD17347345CD17C3C3FC3010FF4F33310CCF0C00DFF03003;
defparam sp_inst_8.INIT_RAM_16 = 256'h075C307570CFC3F0C00F3CFD0300030D0D18030C358034600D180318030C30C0;
defparam sp_inst_8.INIT_RAM_17 = 256'h30C78C30FF0C004D30C0075C307570CFF075C307570CFC3F0C0075C307570CFF;
defparam sp_inst_8.INIT_RAM_18 = 256'h007C71BC300373F0C00C30CF0C00D4CC34CCD4CC34CC0CD4CCD3334CC35330C5;
defparam sp_inst_8.INIT_RAM_19 = 256'hC00D74C344CFC30030C30C8F0C003330C335D4D4CCD737F7E0CC3E3F03001B0C;
defparam sp_inst_8.INIT_RAM_1A = 256'h0C00D130F3C300CF333C3000F3D47DF147CCCF75C0C00345773FC0C000CF3DC0;
defparam sp_inst_8.INIT_RAM_1B = 256'hF321C804FFD771FDDFFD03003FC7013FF77013FF5DC7CDC04FFD7417FDDFFDD4;
defparam sp_inst_8.INIT_RAM_1C = 256'h703430F0C000C030CCC7FF3C330FF0C033C330C0C3007CFEC0804FFD32013FB5;
defparam sp_inst_8.INIT_RAM_1D = 256'h00530C230CF0C00D0D0340DC340D40D7030F0C0034DC35035030F0C003435C0D;
defparam sp_inst_8.INIT_RAM_1E = 256'h0C00434F034D3DD430010D34F034F750C00330C00330C07F034F4301FC0D3D0C;
defparam sp_inst_8.INIT_RAM_1F = 256'hCF3B1CCCFCCF3CCD77CC0C00CDF0CE7FCCF33E7FCCF27CCCCCD030033CF5DCF4;
defparam sp_inst_8.INIT_RAM_20 = 256'h3C3000CC0CCF0C00C0CCC30C323C3001CCC733134C31CCC330CC33C3002C7C43;
defparam sp_inst_8.INIT_RAM_21 = 256'hC3330CC3330CC33DC30001701D030010D0C7CF0C07CC1CFC30017D30CC134C33;
defparam sp_inst_8.INIT_RAM_22 = 256'h1030CC6150340340341740D0F335440D337140D0CDC030FC0C04F0C00C3330CC;
defparam sp_inst_8.INIT_RAM_23 = 256'h10FF003CD1F3FC00F343AFF003CD3D3FC00F38FF003C0380C0141818141030D4;
defparam sp_inst_8.INIT_RAM_24 = 256'h03030FC0C017FCCC50F313C33D10CC0F10C000C3F030143D1FF003C43FC00F14;
defparam sp_inst_8.INIT_RAM_25 = 256'h30053F10F10C080FC0C014FD10F10C080FC0C017FCC8434C84D30CF443303C43;
defparam sp_inst_8.INIT_RAM_26 = 256'h1F0FCCC0F3FCCC30C0F3FC30CF3FC30CF3FC30C0C30F0F333300CCC00C0303F0;
defparam sp_inst_8.INIT_RAM_27 = 256'h5DF3B2803005CF3F35034C0D33F3C43F10FC4FC03005F2F3CBD0FD0C3C0FC0C0;
defparam sp_inst_8.INIT_RAM_28 = 256'hF397CC3D90E41910CE905434684337D90E80A031A10FC0C0173CE85DF3A33CEC;
defparam sp_inst_8.INIT_RAM_29 = 256'hCF3DF90F90F90C24DD0E4F03005082038543450432905434544309097F6430CC;
defparam sp_inst_8.INIT_RAM_2A = 256'h73F03005707370C7370C7370F50F50C1C0FC0C0177CF50C10C343F03005DFE3F;
defparam sp_inst_8.INIT_RAM_2B = 256'hD0F1D3CF346031170D586186045C3FF00C63C03004CD80C3D03005AF50C1C90E;
defparam sp_inst_8.INIT_RAM_2C = 256'hF7DF7000F4030C30C330CC3C743C743C743C743C743C74F1D0F1D0F1D0F1D0F1;
defparam sp_inst_8.INIT_RAM_2D = 256'hC330CC3C643C643C643C643C643C64F190F190F190F193CF303031170C17DF7D;
defparam sp_inst_8.INIT_RAM_2E = 256'hF0300170FF0FFFFFFFF1F40C73DC34150CD13F431D70C77DF7DF70E0F4030C30;
defparam sp_inst_8.INIT_RAM_2F = 256'hC2C0FC0C0155FF1FC7C4C3DD0F743DD0F80C03F03004375FC0C014FD0C3003C3;
defparam sp_inst_8.INIT_RAM_30 = 256'hFA177C3130C33300C28A283D90F4030C30F90F90FC0C01687D5F73F733F90F90;
defparam sp_inst_8.INIT_RAM_31 = 256'hF033333030050308005CC7B305CC7B307B30330C31333E430903F030051F30FF;
defparam sp_inst_8.INIT_RAM_32 = 256'h0C014182C32C3D430703F03005FF3F3CDC03CCF3FFCC4DCFCF30D3CF0D0C4DCC;
defparam sp_inst_8.INIT_RAM_33 = 256'hCF80F50C140FC0C0154FF31D3D4CF310F4CF3CCF94F50C180FC0C01187D030FC;
defparam sp_inst_8.INIT_RAM_34 = 256'hD0FC87DC30FFC0C01743F3310C0C0FC0C014CFF3033CC014CF43C433C3CC74FC;
defparam sp_inst_8.INIT_RAM_35 = 256'h310300513FCC4CF304533D0F10CF0F3DD3F33E208FF32374FCF310F4CF3CCF8C;
defparam sp_inst_8.INIT_RAM_36 = 256'h1433CFCD43C0C0F033CF30434F3CF3033C3C0C05FC3005FC0C01037CCCC174C5;
defparam sp_inst_8.INIT_RAM_37 = 256'h24000C000CE0003000338000C000CE0003000338000C000CF040300033C100C0;
defparam sp_inst_8.INIT_RAM_38 = 256'h80300332C200C00CC80C03000320300C000E80C03000364300C000C90C030003;
defparam sp_inst_8.INIT_RAM_39 = 256'hC00CC50403003328100C00CCA0403003328200C00CCB080300332C200C00CCB0;
defparam sp_inst_8.INIT_RAM_3A = 256'h239C000C008D40003003310000C00CC40003003310000C00CC50403003314100;
defparam sp_inst_8.INIT_RAM_3B = 256'h337F0F0D4200C0C008C60C03002318300C008C60C0300231C300C008C70C0300;
defparam sp_inst_8.INIT_RAM_3C = 256'h003000430C430F10C0C030C0C3000070303C43FD0C0C00B0C0C0C00CF300E01F;
defparam sp_inst_8.INIT_RAM_3D = 256'h000000000000000006420013103000CC0E7CC30331F30CC9190F0C0C0001F30C;
defparam sp_inst_8.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3F = 256'hC3F4D01314404C402226FC0001100920841C44410C4D404EF010C801C3410000;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[29:0],sp_inst_9_dout[21:20]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[21:20]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b01;
defparam sp_inst_9.BIT_WIDTH = 2;
defparam sp_inst_9.BLK_SEL = 3'b000;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000000C008F304F00034001131;
defparam sp_inst_9.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_08 = 256'hFFC0C3C3C3040CFCC1500B0C3C30FFFFFFFFFC2022222220000023FFFFFFFFF0;
defparam sp_inst_9.INIT_RAM_09 = 256'h3003F3CF77F77DCCC1F3CFFF70C00FFFFFFFFFFFFFFFCF030FC3FFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_0A = 256'h3FCC87FC8C3FCF30DF21FF230F3CC37CFC30021FFC8CF7F321FCF233FCC37CFC;
defparam sp_inst_9.INIT_RAM_0B = 256'h03004FD3D3FFF03003D3FCC0C00C700C01FD3F30300238C8E30C009F8C8E30C0;
defparam sp_inst_9.INIT_RAM_0C = 256'hC0037D03003FF4FEF3EF3EF3FC0C00FFF4FFBCFBCFBCFF03003F4FFBCFBCFBFF;
defparam sp_inst_9.INIT_RAM_0D = 256'h0000C0C017F3CF7C0CC0C017FFD8B22C3D37F3CD57FFCF8BF7C8BCFCCDCCFFC0;
defparam sp_inst_9.INIT_RAM_0E = 256'hCF0CF3DC4CCF3DC4CCF3DC4CCF3DC0CCF3DC4CCF3D8CCF3D30700C73C0F1F3FF;
defparam sp_inst_9.INIT_RAM_0F = 256'h33388CC33CE78C3FC3005C7F3DF030CF073C1CF3DC734CFC1CF073CF71CD33CC;
defparam sp_inst_9.INIT_RAM_10 = 256'h303D0C00730C030CCF7703F33C30003C30000C000C00030000C00FC8CDC300CC;
defparam sp_inst_9.INIT_RAM_11 = 256'h005FFF62C8B0F4DFCF355FFF3E2FDF22F3F33733FF03005FCF3DF03303003F03;
defparam sp_inst_9.INIT_RAM_12 = 256'h71333CF71333CF71333CF70333CF71333CF6333CF4C18031CF03C7CFFC000303;
defparam sp_inst_9.INIT_RAM_13 = 256'h0C0171FCFFC00E088CF7C0C33C1CF073CF71CD33F073C1CF3DC734CF333C33CF;
defparam sp_inst_9.INIT_RAM_14 = 256'h5CF030034F03003FFDCDFFF03005373F1330CCDF03000DCCF030000C000301F3;
defparam sp_inst_9.INIT_RAM_15 = 256'hC30C0F0C00E23388CE2338B388CE23C3C3FC3014FF4F33310CCF0C00D4F03003;
defparam sp_inst_9.INIT_RAM_16 = 256'h075C307570CFC3F0C00F3CFD0300030D0D28830C368834A20D288328831C30C0;
defparam sp_inst_9.INIT_RAM_17 = 256'h30C7CC30FF0C008E30C0075C307570CFF075C307570CFC3F0C0075C307570CFF;
defparam sp_inst_9.INIT_RAM_18 = 256'h007C713C300373F0C00C30CF0C00D4CC34CCD4CC34CC0CD4CCD3334CC35330C4;
defparam sp_inst_9.INIT_RAM_19 = 256'hC00E78C388CFC30030C30C4F0C003330C339E4E4CCE33BF3E2CC3C3F0300130C;
defparam sp_inst_9.INIT_RAM_1A = 256'h0C00E230F3C300CF333C3000F3E87DF287CCCF75C0C00389BB3FC0C000CF3DC0;
defparam sp_inst_9.INIT_RAM_1B = 256'hF391E408FFD791FE8F7D03003FC9023FF79023FF6E47CE408FFD7A17FE8F7DD4;
defparam sp_inst_9.INIT_RAM_1C = 256'h703430F0C000C030CCC7FF3C330FF0C033C330C0C3007CFFC2408FFD39023FF6;
defparam sp_inst_9.INIT_RAM_1D = 256'h00730C030CF0C00D0D0340D0360D40D7030F0C0034DC35035030F0C003435C0D;
defparam sp_inst_9.INIT_RAM_1E = 256'h0C00534F134D3DD430014D34F134F750C00330C00330C06E134F4301B84D3D0C;
defparam sp_inst_9.INIT_RAM_1F = 256'hCF371DCCDCCF3DCD76CC0C00CDF0CF7FCCF33F7FCCF37CCCCCD030033CF5ECF4;
defparam sp_inst_9.INIT_RAM_20 = 256'h3C3000CC0CCF0C00C8CCC30C303C3001CCC733238C31CCC330CC33C3001C7C83;
defparam sp_inst_9.INIT_RAM_21 = 256'hC3330CC3330CD33DC3000C70CD030020E0C7CF0C07CC1CFC30027E30CC238C33;
defparam sp_inst_9.INIT_RAM_22 = 256'h113CCC71513C13C13C1B44F0F336C44F337144F0CDC030FC0C04F0C00C3330CC;
defparam sp_inst_9.INIT_RAM_23 = 256'h20FF003871F3FC00E1C30FF003873F3FC00E1CFF003C0340C0141C1C1B113CDB;
defparam sp_inst_9.INIT_RAM_24 = 256'h06030FC0C017FCD861F617C33D10CC0F10C1C0C3F030143E1FF003C83FC00F28;
defparam sp_inst_9.INIT_RAM_25 = 256'h30053F10F10C180FC0C014FD10F10C180FC0C017FCD8474D85D30CF443303C43;
defparam sp_inst_9.INIT_RAM_26 = 256'h1F1FCC20F77CCC3020F77C30CF77C30CF77C30C0C30F1F333300CCC00C0303F0;
defparam sp_inst_9.INIT_RAM_27 = 256'h59B310403005CF3135134C4D3310443110C44C40300512F04BD0FD0C040FC0C0;
defparam sp_inst_9.INIT_RAM_28 = 256'hF397CC3DD0C41510CA109838544327DD0C401031510FC0C0173CC459B3133CC4;
defparam sp_inst_9.INIT_RAM_29 = 256'hCF39FD0FD0FD0C04990C4F0300501043C983854432109838544301097F7430CC;
defparam sp_inst_9.INIT_RAM_2A = 256'h03F03005000370C0370C0370FD0FD0C000FC0C01450FD0C040313F030059F43D;
defparam sp_inst_9.INIT_RAM_2B = 256'hD0D1D3CF300031570C400000055C3FF00003C03004CC00C3D03005CFD0C0010C;
defparam sp_inst_9.INIT_RAM_2C = 256'hFBEFB000F4030C30C330CC3D7434743D7434743D743474F5D0D1D0F5D0D1D0F5;
defparam sp_inst_9.INIT_RAM_2D = 256'hC330CC3D7434743D7434743D743474F5D0D1D0F5D0D1D3CF303031570C57EFBE;
defparam sp_inst_9.INIT_RAM_2E = 256'hF030017CFFCFFFFFFFC1FC0C73CC3C2610E53E431170C7BEFBEFB0F0F4030C30;
defparam sp_inst_9.INIT_RAM_2F = 256'hC380FC0C0155FE1F87C4C3D90F643D90F80F03F03004775FC0C015F90C3C43F3;
defparam sp_inst_9.INIT_RAM_30 = 256'hFE11FC3030C73300C38E383D90F4030C30F90F90FC0C01787D5F62E722F90F90;
defparam sp_inst_9.INIT_RAM_31 = 256'hF03333303005230E004CC7F304CC7F307F30330C31333E430E03F030051F30FF;
defparam sp_inst_9.INIT_RAM_32 = 256'h0C014343C33C3E430D03F03005FF3F3CF407CCF3FFCC4DCFCF30D7CF0F804DCC;
defparam sp_inst_9.INIT_RAM_33 = 256'hCF34F90C340FC0C0174FF3DC7F4CF321F5DF3CCF34F90C340FC0C01347DC30FC;
defparam sp_inst_9.INIT_RAM_34 = 256'h94EF07D830FFC0C01653BC390C300FC0C0170FF3D33CCD15DF47C877C7CF71FC;
defparam sp_inst_9.INIT_RAM_35 = 256'h3103005C3FCF0CF330577D1F21DF1F39C7F33CC30FF3C271FCF321F5DF3CCF30;
defparam sp_inst_9.INIT_RAM_36 = 256'h1433CECD47C4C1F133CF30535F3CF313383C0C05FC3005FC0C01037CCCC078C6;
defparam sp_inst_9.INIT_RAM_37 = 256'h2C000C000CB000300032C000C000CB000300032C000C000CB000300032C000C0;
defparam sp_inst_9.INIT_RAM_38 = 256'hC03003328300C00CEB0C0300036C300C000CB0C0300032C300C000CB0C030003;
defparam sp_inst_9.INIT_RAM_39 = 256'hC00CCA0C03003328300C00CCA0C03003328300C00CCA0C03003328300C00CCA0;
defparam sp_inst_9.INIT_RAM_3A = 256'h3324300C00CCA0C03003328300C00CCA0C03003328300C00CCA0C03003328300;
defparam sp_inst_9.INIT_RAM_3B = 256'h337F0F0E4200C0C00CC90803003324200C00CC908030033A4200C00CD9080300;
defparam sp_inst_9.INIT_RAM_3C = 256'h403901430C430F00C0C030C0C3002470303C83F80C0C00F0C0C0C00CF304D01F;
defparam sp_inst_9.INIT_RAM_3D = 256'h00000000000000000BFA0028203000CC0C7CC30381F30E00100F0C0C0001F30E;
defparam sp_inst_9.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3F = 256'hA3B8ABA2ACAE8AB0323BA8CC9310F3CF0C00408E28B7A38AA3BBCA3EA0BA8000;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[29:0],sp_inst_10_dout[23:22]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[23:22]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b01;
defparam sp_inst_10.BIT_WIDTH = 2;
defparam sp_inst_10.BLK_SEL = 3'b000;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000011822CB2003A2232228880;
defparam sp_inst_10.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_08 = 256'hAA80D1E1D100AEE9E002AEE81D14AAAAAAAAA81111111111111112AAAAAAAAA0;
defparam sp_inst_10.INIT_RAM_09 = 256'hA29AB82222A228A90410AAA62A808AAAAAAAAAAAAAAA8EDB658AAAAAAAAAAAAA;
defparam sp_inst_10.INIT_RAM_0A = 256'h7AA8429D453AAAA04A10A7514BAA8128AAA2910A9D45E2AA10A4B517AA8128AA;
defparam sp_inst_10.INIT_RAM_0B = 256'hAA2A1BCACAC02AA2A7CAF2AA8A9D36A8A83CACAAA291944651A8A44944651A8A;
defparam sp_inst_10.INIT_RAM_0C = 256'h8A9100AA2A7EB2B1A61A618AAAA8A9FEB2BC69869862AAAA2A7F2BC69869862A;
defparam sp_inst_10.INIT_RAM_0D = 256'hAAAAAA8A8302AB0E20AA8A83AAC66198A802A28802AEAA02828028A8E888AAAA;
defparam sp_inst_10.INIT_RAM_0E = 256'hAB8AAACA28AAACA28AAACA28AAACAA8AAACA28AAAC68AAACA221282AA200A2AA;
defparam sp_inst_10.INIT_RAM_0F = 256'hA225488A289248A8AA2A0C2AAC3881EF82AE0AAA882A28BE0AB82AAA20A8A2A8;
defparam sp_inst_10.INIT_RAM_10 = 256'h4290A8A629A4A9A6A62229A62AA2922AA292A8A4A8A4AA292A8A42D490AA2908;
defparam sp_inst_10.INIT_RAM_11 = 256'h2A0EAB198662A00A8A200ABAA80A0A00A2A3A222AAAA2A0C0AAC3882AA298790;
defparam sp_inst_10.INIT_RAM_12 = 256'h28A2AAB28A2AAB28A2AAB2AA2AAB28A2AAB1A2AAB28884A0AA88028AAAAAAAAA;
defparam sp_inst_10.INIT_RAM_13 = 256'hA8A830AABA954A0028B0E207BE0AB82AAA20A8A2F82AE0AAA882A28AA2AE2AAB;
defparam sp_inst_10.INIT_RAM_14 = 256'h08AAA2A71AAA2A7EAC8CBAAAA2A0A2AA0AA2AA8EAA2A68EAAAA292A8A4AA28A2;
defparam sp_inst_10.INIT_RAM_15 = 256'h8A088AA8A495625589562562558956A9A9AAA280AA0B2A200A8AA8A9C2AAA2A7;
defparam sp_inst_10.INIT_RAM_16 = 256'h210A92102A4A8AAA8A9E3808AA2989A44850224A91022140885022502284A088;
defparam sp_inst_10.INIT_RAM_17 = 256'h9A62E692AAA8A4651A8A610A92102A4AA210A92102A4A8AAA8A610A92102A4AA;
defparam sp_inst_10.INIT_RAM_18 = 256'hA6252A5AA29A2AAA8A6AAAAAA8A682A8A2AA82A8A2A8AA82AA8AAA2A8A0AA2A0;
defparam sp_inst_10.INIT_RAM_19 = 256'h8A492482648AAA29228A2A8AA8A9122282249090889626A680A8AA2AAA29A5A8;
defparam sp_inst_10.INIT_RAM_1A = 256'hA8A4992102AA29D0202AA2A490B8008380200800AA8A9264662AAA8A924220AA;
defparam sp_inst_10.INIT_RAM_1B = 256'h55E078047740E0095554AA2A776E011DD0E011DD1781578047740E0009555042;
defparam sp_inst_10.INIT_RAM_1C = 256'h212124AA8A6A4A92AA6227AA92A6AA8A7AA92A626A2A00776B8047748E011DD1;
defparam sp_inst_10.INIT_RAM_1D = 256'hA629A4A9A4AA8A644852148521480482125AA8A6908520120124AA8A69120848;
defparam sp_inst_10.INIT_RAM_1E = 256'hA8A6091189104002A29824411891000A8A699A8A699A8A1589152A28562454A8;
defparam sp_inst_10.INIT_RAM_1F = 256'hEAAE0898B8EAA898318AA8A9EC365F2022089B22220B2222220AA2A796701442;
defparam sp_inst_10.INIT_RAM_20 = 256'h2AA29964A64AA8A6A8A8AAAAAA2AA2986A61A91944A86A6A9AA699AA2A780169;
defparam sp_inst_10.INIT_RAM_21 = 256'h8AAAAA8AAAA80AA0AA2A4B0AB0AA291A526266A8A28A0A6AA291251964194699;
defparam sp_inst_10.INIT_RAM_22 = 256'h0868A8E008688688680E21A0AA33821A2AE021A28B80A2AAA8A1AA8A68AAAAAA;
defparam sp_inst_10.INIT_RAM_23 = 256'hBAEA5528E0ABA954A38AAEA5528E2A3A954A38EA5528A9EA8A8138380E0868CE;
defparam sp_inst_10.INIT_RAM_24 = 256'h2E0A2AAA8A83AAB810AE0286280A8A2A0A8B828AAAA282AF8EA5528EBA954A3E;
defparam sp_inst_10.INIT_RAM_25 = 256'hA2A0AA0AA0A8B82AAA8A80200AA0A8B82AAA8A83AAB8221B808618A02A28A82A;
defparam sp_inst_10.INIT_RAM_26 = 256'h8B0AA9E0A228A8A0E0A228A28A228A28A228A2828A2A0A2A2A888AA2288A22AA;
defparam sp_inst_10.INIT_RAM_27 = 256'h0C62E38AA2A0EAAE20891A2462E3829E0A78278AA2A0E3AB8ECAACA8B82AAA8A;
defparam sp_inst_10.INIT_RAM_28 = 256'h08C000A0CAB80E0A8FE045E5382A300CAB82E0A0E0AAAA8A83AAB80C62E3AAB8;
defparam sp_inst_10.INIT_RAM_29 = 256'h8A6CACAACAACA8B8CC2B8AAA2A02E383C45E5382A3E045E5382A2E0C0032A28E;
defparam sp_inst_10.INIT_RAM_2A = 256'hE2AAA2A0E0E2E28E2E28E2E2ACAACA8B82AAA8A8308ACA8B8CAE2AAA2A0CA228;
defparam sp_inst_10.INIT_RAM_2B = 256'hC288C2AAA2E0A0C2A838E38E030AAAAAA8E2AAA2A10B82080AA2A0BACA8B8C2B;
defparam sp_inst_10.INIT_RAM_2C = 256'h861862E0A08A28A28A2288A830A230A830A230A830A230A0C288C2A0C288C2A0;
defparam sp_inst_10.INIT_RAM_2D = 256'h8A2288A830A230A830A230A830A230A0C288C2A0C288C2AAA2E0A0C2A8C21861;
defparam sp_inst_10.INIT_RAM_2E = 256'hAAA2A828AA8AA2222238A8282698A811C8922B2A0C2A8061861862A0A08A28A2;
defparam sp_inst_10.INIT_RAM_2F = 256'h8A82AAA8A8304A068040040CA832A0CAA82A0AAAA2A1D2CAAA8A83ACA8A8CAA2;
defparam sp_inst_10.INIT_RAM_30 = 256'hAA04AA9A9A6296224A8A2828CAA08A28A2ACAACAAAA8A82800C5159215ACAACA;
defparam sp_inst_10.INIT_RAM_31 = 256'h9A9A9A9AA2A0A92A060662D920662D922D90A228A8192B2A2A0AAAA2A08B9A7A;
defparam sp_inst_10.INIT_RAM_32 = 256'hA8A80A824A24AB2A2A0AAAA2A0DAAEAAA823A8A276AA348BAAAA838AA68E1488;
defparam sp_inst_10.INIT_RAM_33 = 256'h8AA8ACA8A82AAA8A828EAA8A2A8EAA10A04A298AA8ACA8A82AAA8A868148926A;
defparam sp_inst_10.INIT_RAM_34 = 256'h80AA8148926AAA8A8202AA2CA8A82AAA8A828EAAA3AA8A004A028412828A28A9;
defparam sp_inst_10.INIT_RAM_35 = 256'h98AA2A0A3AAA8EAA2801280A104A0A28A2A62AA28EAAA228AEAA10A04A298AA8;
defparam sp_inst_10.INIT_RAM_36 = 256'h8032AA8821A0886822CAAA02062CAA822A2AA8A0AAA2A0EAA8A8792AAAA32A62;
defparam sp_inst_10.INIT_RAM_37 = 256'hA8A2A8A9E6A28AA2A79A8A2A8A9E6A28AA2A79A8A2A8A9E6A28AA2A79A8A2A8A;
defparam sp_inst_10.INIT_RAM_38 = 256'h8AA2A6928A2A8A9A6A28AA2A79A8A2A8A9E6A28AA2A79A8A2A8A9E6A28AA2A79;
defparam sp_inst_10.INIT_RAM_39 = 256'h8A9A4A28AA2A6928A2A8A9A4A28AA2A6928A2A8A9A4A28AA2A6928A2A8A9A4A2;
defparam sp_inst_10.INIT_RAM_3A = 256'h6928A2A8A9A4A28AA2A6928A2A8A9A4A28AA2A6928A2A8A9A4A28AA2A6928A2A;
defparam sp_inst_10.INIT_RAM_3B = 256'h262AA6A68A226A8A9A4A28AA2A69A8A2A8A9A5A28AA2A6928A2A8A9A4A28AA2A;
defparam sp_inst_10.INIT_RAM_3C = 256'h829A08862A09A65A6A8A42626A2A681A98916955A6A8A9AA626A8A9EAA21A04A;
defparam sp_inst_10.INIT_RAM_3D = 256'h000000000000000004012A6A2AA2A4A4A7004429A001128E0E1026A8A948B9A6;
defparam sp_inst_10.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3F = 256'h5044511110444440111514005014000005144441141540414010140140110000;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[29:0],sp_inst_11_dout[25:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[25:24]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b01;
defparam sp_inst_11.BIT_WIDTH = 2;
defparam sp_inst_11.BLK_SEL = 3'b000;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000020D330D3003937737640C0;
defparam sp_inst_11.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_08 = 256'h5550F9E5F9208FE8F803F4185F98000000000103000000333333315555555554;
defparam sp_inst_11.INIT_RAM_09 = 256'h62343A69001004248CA141551980C0000000000000001C27C449555555555555;
defparam sp_inst_11.INIT_RAM_0A = 256'hF061201F27306186404807C9C7861900566234821F27C21848047C9F06190056;
defparam sp_inst_11.INIT_RAM_0B = 256'h96202BCACAD569620FCAF665883F3E5880BCAD996234D25349988D0925349988;
defparam sp_inst_11.INIT_RAM_0C = 256'h8831249620FC32B410410419565883FC32BD04104106559620FF2BD041041065;
defparam sp_inst_11.INIT_RAM_0D = 256'h955565880318632E2065880318C2008084028004000C610012000050E4001565;
defparam sp_inst_11.INIT_RAM_0E = 256'h638618C200618C200618C200618C280618C200618C00618C0020280862180146;
defparam sp_inst_11.INIT_RAM_0F = 256'h844321186102218566200C018CB883EF808E02184808207E0238086120208160;
defparam sp_inst_11.INIT_RAM_10 = 256'hD0D4988D2D347D3535030D50066233066233988C988CE6233988D8F234662361;
defparam sp_inst_11.INIT_RAM_11 = 256'h200C63080202100A0010003184004800014390005596200C618CB881962367B2;
defparam sp_inst_11.INIT_RAM_12 = 256'h0801863080186308018630A01863080186300186300080A0218860051A555596;
defparam sp_inst_11.INIT_RAM_13 = 256'h98803006363FC7002032E20FBE02380861202081F808E02184808205818E1863;
defparam sp_inst_11.INIT_RAM_14 = 256'h0C19620F019620FC1C8CB559620000060000010D9620D0D1196233988CE62011;
defparam sp_inst_11.INIT_RAM_15 = 256'h1820A1988D0C043010C043043010C04D4D5662021823180006059883C219620F;
defparam sp_inst_11.INIT_RAM_16 = 256'h1102111008410859883C309496235D74E0002821D0028000A00028002845820A;
defparam sp_inst_11.INIT_RAM_17 = 256'hD35374D015988D349988D102111008418110211100841085988D102111008418;
defparam sp_inst_11.INIT_RAM_18 = 256'h8D0407566234005988D18611988D000040010000400081000100040004000010;
defparam sp_inst_11.INIT_RAM_19 = 256'h88D0220432016623461861C19883148608408202210040604001871596237598;
defparam sp_inst_11.INIT_RAM_1A = 256'h588D0C83986623F98186620D963824A382788110658834300005658836580465;
defparam sp_inst_11.INIT_RAM_1B = 256'h9EE0B8027742E09809E49620F76E009DD2E009DD0B827B8027742E029809E442;
defparam sp_inst_11.INIT_RAM_1C = 256'h3080821988DB46D213530784D1355988F84D1357662026776B802774AE009DD0;
defparam sp_inst_11.INIT_RAM_1D = 256'h8D2D347D341988D4E0C8320C832002030821988DD20C800800821988DD380C20;
defparam sp_inst_11.INIT_RAM_1E = 256'h588D0D0B0D08244262343420B0D0910988DD1988DD19880C0D09262030342498;
defparam sp_inst_11.INIT_RAM_1F = 256'hE18E008078E1848030065883ECBC7F2566599F26665B26666649620FA6B08852;
defparam sp_inst_11.INIT_RAM_20 = 256'h066237447441988D1C1C1861870662344051014D24044050D435D56620F8270D;
defparam sp_inst_11.INIT_RAM_21 = 256'h00048100048180046620C8268496234F4B5045988046005662342497444D25D1;
defparam sp_inst_11.INIT_RAM_22 = 256'h000860E000080080080C00205033800218E000220780821658835988D0004810;
defparam sp_inst_11.INIT_RAM_23 = 256'hBAD8FF1CE01B63FC7389CD8FF1CE06363FC738D8FF1C6DE5880338380E0008CE;
defparam sp_inst_11.INIT_RAM_24 = 256'h2E08216588030638080E000C14020621020B82085962026F8D8FF1CEB63FC73E;
defparam sp_inst_11.INIT_RAM_25 = 256'h620041021020B82165880184021020B821658803063800038000305008188408;
defparam sp_inst_11.INIT_RAM_26 = 256'h038063E060002080E0600082060008206000820208218019198A0662A0A82859;
defparam sp_inst_11.INIT_RAM_27 = 256'h0C01E3896200E18E000D003401E380DE037807896200E30B8DC21C20B8216588;
defparam sp_inst_11.INIT_RAM_28 = 256'h9AC28484C2380E020FE002C23808324C2382E080E02165880386380C01E38638;
defparam sp_inst_11.INIT_RAM_29 = 256'hC10C9C21C21C20B8CC2385962002E383C02C238083E002C238082E0C2930820E;
defparam sp_inst_11.INIT_RAM_2A = 256'hE0596200E0E0C20E0C20E0C21C21C20B8216588030C1C20B8C8E0596200C9304;
defparam sp_inst_11.INIT_RAM_2B = 256'hCA08C84102E080C02038E38E0300855008E16562038B828A496200F1C20B8C23;
defparam sp_inst_11.INIT_RAM_2C = 256'h104102E01088208208020084328232843282328432823210CA08CA10CA08CA10;
defparam sp_inst_11.INIT_RAM_2D = 256'h08020084328232843282328432823210CA08CA10CA08C84102E080C020C24104;
defparam sp_inst_11.INIT_RAM_2E = 256'h596200380380199999B8B8201C40B800CC0307080C020104104102E010882082;
defparam sp_inst_11.INIT_RAM_2F = 256'h0B8216588030AE0B8240824C213084C2382E08596203D2C96588031C20B8C8E0;
defparam sp_inst_11.INIT_RAM_30 = 256'h8E00C4D7D350D0134B8E3804C2108820821C21C21658803824C90C03001C21C2;
defparam sp_inst_11.INIT_RAM_31 = 256'h56D6D6D962007D2E0D0453511045351135108020841107082E085962004DD371;
defparam sp_inst_11.INIT_RAM_32 = 256'h58800B83483487082E08596200D18C8638010041746114C321840104478D14C0;
defparam sp_inst_11.INIT_RAM_33 = 256'h05B85C20B8216588038C18C2038E184800401405B85C20B82165880F824D9656;
defparam sp_inst_11.INIT_RAM_34 = 256'hC033824D965565880300CE1C20B8216588038C18E3860E004020021020070804;
defparam sp_inst_11.INIT_RAM_35 = 256'hD896200E30638E18380100800840801C201016E38C18E3080E184800401405B8;
defparam sp_inst_11.INIT_RAM_36 = 256'h007063800101004041C18404041C18441E165880566200D65880FD2666732F63;
defparam sp_inst_11.INIT_RAM_37 = 256'hB8A25883F6E289620FDB8A25883F6E289620FDB8A25883F6E289620FDB8A2588;
defparam sp_inst_11.INIT_RAM_38 = 256'h89620FD38A25883F7E289620FDB8A25883F6E289620FDB8A25883F6E289620FD;
defparam sp_inst_11.INIT_RAM_39 = 256'h883F4E289620FD38A25883F4E289620FD38A25883F4E289620FD38A25883F4E2;
defparam sp_inst_11.INIT_RAM_3A = 256'hFD38A25883F4E289620FD38A25883F4E289620FD38A25883F4E289620FD38A25;
defparam sp_inst_11.INIT_RAM_3B = 256'h1D0135378A1365883F5E289620FD38A25883F4E289620FD38A25883F4E289620;
defparam sp_inst_11.INIT_RAM_3C = 256'h81DE0080210D35C36588DB536620F826D4D70D70365883D35365883E180020C0;
defparam sp_inst_11.INIT_RAM_3D = 256'h000000000000000005A920FE39620DB5B7264E6DE0993B8E0E39B65883C4DD37;
defparam sp_inst_11.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3F = 256'h51700D5200254800101840001014514503340C003C95200510100C00C2058000;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[29:0],sp_inst_12_dout[27:26]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[27:26]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b01;
defparam sp_inst_12.BIT_WIDTH = 2;
defparam sp_inst_12.BLK_SEL = 3'b000;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'h000000000000000000000000000000000000000000DD14451451728470448810;
defparam sp_inst_12.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_08 = 256'hAA97090909A32400480806E39095AAAAAAAAA91011111144444406AAAAAAAAA5;
defparam sp_inst_12.INIT_RAM_09 = 256'h8C8AB28A22A2288880A2AAAA22351AAAAAAAAAAAAAAA96D82692AAAAAAAAAAAA;
defparam sp_inst_12.INIT_RAM_0A = 256'h2A8A2294242A8A2A4A88A5090B28A928A88C88889424A0A288A48092A8A928A8;
defparam sp_inst_12.INIT_RAM_0B = 256'h28CA2140406A828CA140588A328410A3289406228C8812604923220126049232;
defparam sp_inst_12.INIT_RAM_0C = 256'h32852828CA169018A28A28A2A8A32856901628A28A28AA28CA1501628A28A28A;
defparam sp_inst_12.INIT_RAM_0D = 256'h2AAA8A3281AA8924C88A3280A24020082820228802A68A32A08328A84898AA8A;
defparam sp_inst_12.INIT_RAM_0E = 256'h8908A248288A248288A248288A248288A248288A24288A24AE0C82228CA8A2A8;
defparam sp_inst_12.INIT_RAM_0F = 256'h2AA02AA28A802A2A88CA062A24932041222488A2822208848892228A08882288;
defparam sp_inst_12.INIT_RAM_10 = 256'h2218232201848186862061A2288C84688C842321232108C842322A028888C8AA;
defparam sp_inst_12.INIT_RAM_11 = 256'hCA0289008020A0808A200A9A28CA820CA2A12262AA28CA06AA24932228C8A602;
defparam sp_inst_12.INIT_RAM_12 = 256'h20A228920A228920A228920A228920A22890A22892B832088A32A28AA0AAAA28;
defparam sp_inst_12.INIT_RAM_13 = 256'h232818A89880085308924C81048892228A0888221222488A2822208A22242289;
defparam sp_inst_12.INIT_RAM_14 = 256'h01A28CA10A28CA1AA4041AA28CA0A2A80AAAAA8628CA286AA28C84232108C8A2;
defparam sp_inst_12.INIT_RAM_15 = 256'hA26A2A2322802A00A802A02A00A802A1A1A88C82A22AA2A0688A232840A28CA1;
defparam sp_inst_12.INIT_RAM_16 = 256'h21089210225A82A2328618A828C8918428030A2A1030A00C28030A030A9626A2;
defparam sp_inst_12.INIT_RAM_17 = 256'h18604612AA232204923221089210225A221089210225A82A23221089210225A2;
defparam sp_inst_12.INIT_RAM_18 = 256'h222428588C8A2AA2322A28AA232282A8A2AA82A8A2AB2A82AA8AAA2A8A0AA6A1;
defparam sp_inst_12.INIT_RAM_19 = 256'h3228028A028A88C8A8A28A1A23285AA88AA00282AA82A2828CAA286A28C88523;
defparam sp_inst_12.INIT_RAM_1A = 256'hA32280A0AA88C84AA2A88CA21A93282132889A208A328A00226A8A32886A688A;
defparam sp_inst_12.INIT_RAM_1B = 256'hA24C934255424CA00A2828CA1544D095524D095509328934255424C2A00A2880;
defparam sp_inst_12.INIT_RAM_1C = 256'h04A0A2A23220481CA860672A1286A23232A1286448CA2A554134255424D09550;
defparam sp_inst_12.INIT_RAM_1D = 256'h2201848184A23224280A0280A02812804A2A23221280A04A04A2A232210A0128;
defparam sp_inst_12.INIT_RAM_1E = 256'hA3220108810828808C8804208810A2023221923221923200810A08C802042823;
defparam sp_inst_12.INIT_RAM_1F = 256'h4A24C808934A28081088A3284492450A88A2210888A1088888828CA3289088A0;
defparam sp_inst_12.INIT_RAM_20 = 256'h288C8864864A2322A1A1A28A28688C886A61A98124A86A6A1A861988CA132821;
defparam sp_inst_12.INIT_RAM_21 = 256'h9AAA2A8AAA2A8AA888CA13283828C8804862662322880A688C88049864812619;
defparam sp_inst_12.INIT_RAM_22 = 256'hC823884C082382382346208CAA113208E24C208C893228A8A320A23228AAA2AA;
defparam sp_inst_12.INIT_RAM_23 = 256'h106200214CA18800853216200214E8D8800853620021814A3280131344C82344;
defparam sp_inst_12.INIT_RAM_24 = 256'h04D24A8A3280A89308A4C292284888CA48813492A28C80810620021418800854;
defparam sp_inst_12.INIT_RAM_25 = 256'h8CA0AA48A488138A8A3282A848A488138A8A3280A8932209308248A122232922;
defparam sp_inst_12.INIT_RAM_26 = 256'h898A884C822B8B204C822A2C8822A2C8822A2C88A28A8A222232888C8A22CAA2;
defparam sp_inst_12.INIT_RAM_27 = 256'h04224D328CA04A24E0810A04224D3214C85325328CA04DA13648A488138A8A32;
defparam sp_inst_12.INIT_RAM_28 = 256'hA2428B28489344C8854C00201322128489304E244C8A8A3281289304224D2893;
defparam sp_inst_12.INIT_RAM_29 = 256'h1A24248A48A4881344093A28CA004D3140020132214C0020132204C42A122C8C;
defparam sp_inst_12.INIT_RAM_2A = 256'h4EA28CA04C4E6C84E6C84E6CA48A488130A8A328101A48813424EA28CA042068;
defparam sp_inst_12.INIT_RAM_2B = 256'h48804AAAA04E244288134D34D10A2AAAA34E8A8CA0813CB2828CA05A48813409;
defparam sp_inst_12.INIT_RAM_2C = 256'hA28A204CA0328A28B2288A281220122812201228122012A0488048A0488048A0;
defparam sp_inst_12.INIT_RAM_2D = 256'hB2288A281220122812201228122012A0488048A048804AAAA04E244288408A28;
defparam sp_inst_12.INIT_RAM_2E = 256'hA28CA813A93AAAAAAA901388228813000180692244288228A28A204CA0328A28;
defparam sp_inst_12.INIT_RAM_2F = 256'h8138A8A32810A4C9328082848A1228489304E2A28CA050428A3281A48813424E;
defparam sp_inst_12.INIT_RAM_30 = 256'h24C02A18186212244134D32848A0124A28A48A48A8A32813284A008040A48A48;
defparam sp_inst_12.INIT_RAM_31 = 256'h981818128CA08104C2166059216605920592228A2859692204E2A28CA081185A;
defparam sp_inst_12.INIT_RAM_32 = 256'hA32801317217292204E2A28CA09A262893A1A8A2668A14198A2A818A95361418;
defparam sp_inst_12.INIT_RAM_33 = 256'h8A13A488138A8A32813AA248293CA288A04A288A13A488138A8A328132861868;
defparam sp_inst_12.INIT_RAM_34 = 256'h41993286186A8A32810664E488138A8A32813AA24F2884C04A22A212A28920A8;
defparam sp_inst_12.INIT_RAM_35 = 256'h1028CA04EA893CA21301288A884A8A2482A2284D3AA24D20ACA288A04A288A13;
defparam sp_inst_12.INIT_RAM_36 = 256'h8366893821A1A868629A2A060629A28624E8A320A88CA068A328110888850441;
defparam sp_inst_12.INIT_RAM_37 = 256'h130CA328444C328CA11130CA328444C328CA11130CA328444C328CA11130CA32;
defparam sp_inst_12.INIT_RAM_38 = 256'h328CA11530CA328444C328CA11130CA328444C328CA11130CA328444C328CA11;
defparam sp_inst_12.INIT_RAM_39 = 256'h328454C328CA11530CA328454C328CA11530CA328454C328CA11530CA328454C;
defparam sp_inst_12.INIT_RAM_3A = 256'h11530CA328454C328CA11530CA328454C328CA11530CA328454C328CA11530CA;
defparam sp_inst_12.INIT_RAM_3B = 256'h222A868530E44A328454C328CA11530CA328454C328CA11530CA328454C328CA;
defparam sp_inst_12.INIT_RAM_3C = 256'h3214F8328A1186084A32286448CA13281918218084A32868644A328CA2E08C0A;
defparam sp_inst_12.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFC449CA14D28CA206052A42814CA90934040A84A328081185;
defparam sp_inst_12.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_12.INIT_RAM_3F = 256'hB30C0513D0044F402119C444D100A24803340C092C32024F3206112912023FFF;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[29:0],sp_inst_13_dout[29:28]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[29:28]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b01;
defparam sp_inst_13.BIT_WIDTH = 2;
defparam sp_inst_13.BLK_SEL = 3'b000;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000110041040524450448814;
defparam sp_inst_13.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_08 = 256'hAA90094909602440480406609090AAAAAAAAA95055555500000002AAAAAAAAA4;
defparam sp_inst_13.INIT_RAM_09 = 256'h808AA28A22A2288880A6AAAA22000AAAAAAAAAAAAAAA96482782AAAAAAAAAAAA;
defparam sp_inst_13.INIT_RAM_0A = 256'h2A8A2290246A8A2A4A88A4091A28A929A88088889024A0A288A58092A8A929A8;
defparam sp_inst_13.INIT_RAM_0B = 256'h280A2140406A8280A140588A028010A028940622808812604920220126049202;
defparam sp_inst_13.INIT_RAM_0C = 256'h028528280A169018A28A28A2A8A02856901628A28A28AA280A1501628A28A28A;
defparam sp_inst_13.INIT_RAM_0D = 256'h2AAA8A0280AA8924498A0282A240240A28602A9802A28A12A08129A948A8AA8A;
defparam sp_inst_13.INIT_RAM_0E = 256'h8918A248298A248298A248298A248298A248298A24298A24A204822284A8A6A8;
defparam sp_inst_13.INIT_RAM_0F = 256'h2AA02AA28A802A2A880A022A24912446222888A28222099888A2228A08882689;
defparam sp_inst_13.INIT_RAM_10 = 256'h2218202201858186862061A228808028808020202020080802022A02888808AA;
defparam sp_inst_13.INIT_RAM_11 = 256'h0A0A89009028A180AA600A8A284A8204A6A522A2AA280A02AA2491262808A502;
defparam sp_inst_13.INIT_RAM_12 = 256'h20A628920A628920A628920A628920A62890A628928812088A12A29AA0AAAA28;
defparam sp_inst_13.INIT_RAM_13 = 256'h202808A888801841089244911888A2228A0888266222888A2822209A26246289;
defparam sp_inst_13.INIT_RAM_14 = 256'h01A280A10A280A1AA4141AA280A0A2A84AAAAA86280A286AA2808020200808A2;
defparam sp_inst_13.INIT_RAM_15 = 256'hA22A2A2022802A00A802A02A00A802A1A1A88082A229A2A4289A202840A280A1;
defparam sp_inst_13.INIT_RAM_16 = 256'h61089610224AA2A2028658A82808918428010A2A1010A00428010A010A9622A2;
defparam sp_inst_13.INIT_RAM_17 = 256'h18604612AA202204920221089610224A261089610224AA2A20221089610224A2;
defparam sp_inst_13.INIT_RAM_18 = 256'h22242858808A2AA2022A28AA202282A9A2AA82A9A2A92A82AA8AAA2A9A0AA2A1;
defparam sp_inst_13.INIT_RAM_19 = 256'h0228029A028A8808A8A28A1A20285AA88AA00282AA82A28284AA286A28088520;
defparam sp_inst_13.INIT_RAM_1A = 256'hA02280A0AA88080AA6A880A21A91282512889A208A028A00226A8A02886A688A;
defparam sp_inst_13.INIT_RAM_1B = 256'hA2449182554244A00A28280A15446095524609550912891825542442A00A2880;
defparam sp_inst_13.INIT_RAM_1C = 256'h04A0A2A202205814A860652A1686A20212A16864480A2A554118255424609550;
defparam sp_inst_13.INIT_RAM_1D = 256'h2201858184A20224280A0280A02812804A2A20221280A04A04A2A202210A0128;
defparam sp_inst_13.INIT_RAM_1E = 256'hA022010881082880808804208810A2020221920221920200810A080802042820;
defparam sp_inst_13.INIT_RAM_1F = 256'h8A244809918A28081098A0284482450A88A2210888A10888888280A2289089A0;
defparam sp_inst_13.INIT_RAM_20 = 256'h28808865864A2022A1A1A28A286880886A61A98124A86A6A1A8619880A112821;
defparam sp_inst_13.INIT_RAM_21 = 256'hAAAA2AAAAA2A8AA8880A1128182808804862662022980A688088049865812619;
defparam sp_inst_13.INIT_RAM_22 = 256'h482189440821821821062085AA41120862442084991524A8A020A2022AAAA2AA;
defparam sp_inst_13.INIT_RAM_23 = 256'h1022006144A088018512122006146848801851220061814A0280515104482104;
defparam sp_inst_13.INIT_RAM_24 = 256'h44628A8A0282A89108A442826848984A489118A2A28080850220061408801854;
defparam sp_inst_13.INIT_RAM_25 = 256'h80A0AA48A489114A8A0282A848A489114A8A0282A8912209108209A122612922;
defparam sp_inst_13.INIT_RAM_26 = 256'h888A8845822A8A2545822A289822A289822A2894924A8A626212988489224AA2;
defparam sp_inst_13.INIT_RAM_27 = 256'h0426451280A08A2460810A04264512144851251280A045A11648A489114A8A02;
defparam sp_inst_13.INIT_RAM_28 = 256'hA242992848910448954400201122528489144520448A8A028228910426462891;
defparam sp_inst_13.INIT_RAM_29 = 256'h1A24248A48A4891144891A280A0445154002011225440020112244542A122498;
defparam sp_inst_13.INIT_RAM_2A = 256'h46A280A04546649466494664A48A489118A8A028101A489116246A280A042068;
defparam sp_inst_13.INIT_RAM_2B = 256'h48804AAAA445204289114514410A2AAAA1468A80A09118A28280A05A48911489;
defparam sp_inst_13.INIT_RAM_2C = 256'hA28A2444A1228A2892288A281220122812201228122012A0488048A0488048A0;
defparam sp_inst_13.INIT_RAM_2D = 256'h92288A281220122812201228122012A0488048A048804AAAA445204289408A28;
defparam sp_inst_13.INIT_RAM_2E = 256'hA280A811A91AAAAAAA901149228911000180692204289228A28A2444A1228A28;
defparam sp_inst_13.INIT_RAM_2F = 256'h9114A8A02810A449128082848A122848914452A280A050428A0281A489116246;
defparam sp_inst_13.INIT_RAM_30 = 256'h24402A18186212645114512848A1228A28A48A48A8A02811284A008040A48A48;
defparam sp_inst_13.INIT_RAM_31 = 256'h9818181280A0814452166059616605960595224A285929224452A280A081184A;
defparam sp_inst_13.INIT_RAM_32 = 256'hA0281115525529224452A280A09A2A289161A9A6668A141A8A2A819A95161419;
defparam sp_inst_13.INIT_RAM_33 = 256'h9A11A489114A8A02811AA2482918A288A04A689A11A489114A8A028112861868;
defparam sp_inst_13.INIT_RAM_34 = 256'h41991286186A8A028106646489114A8A02811AA2462894404A229212A29920A8;
defparam sp_inst_13.INIT_RAM_35 = 256'h10280A046A8918A25101288A484A8A6482A268451AA24520A8A288A04A689A11;
defparam sp_inst_13.INIT_RAM_36 = 256'h8066891821A19868669A2A060669A2866468A020A880A068A028110888850441;
defparam sp_inst_13.INIT_RAM_37 = 256'h1104A02844441280A111104A02844441280A111104A02844441280A111104A02;
defparam sp_inst_13.INIT_RAM_38 = 256'h1280A115104A02844441280A111104A02844441280A111104A02844441280A11;
defparam sp_inst_13.INIT_RAM_39 = 256'h02845441280A115104A02845441280A115104A02845441280A115104A0284544;
defparam sp_inst_13.INIT_RAM_3A = 256'h115104A02845441280A115104A02845441280A115104A02845441280A115104A;
defparam sp_inst_13.INIT_RAM_3B = 256'h622A868510644A02845441280A115104A02845441280A115104A02845441280A;
defparam sp_inst_13.INIT_RAM_3C = 256'h161448128A1186084A022864480A11281918218084A02868644A0288A220840A;
defparam sp_inst_13.INIT_RAM_3D = 256'h55555555555555554AF20A145280A206052A428144A90914040A84A028181185;
defparam sp_inst_13.INIT_RAM_3E = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sp_inst_13.INIT_RAM_3F = 256'hA1A8CEB3E82ACFA0232D8C88B2283CF3CA2C480E28F2B38AA3E7E83EF0EAD555;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[29:0],sp_inst_14_dout[31:30]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:30]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b01;
defparam sp_inst_14.BIT_WIDTH = 2;
defparam sp_inst_14.BLK_SEL = 3'b000;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000004500000000104010000004;
defparam sp_inst_14.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_08 = 256'h0001404040410440400400010400000000000054555555444444400000000000;
defparam sp_inst_14.INIT_RAM_09 = 256'h0400100000000000100400000010000000000000000004010000000000000000;
defparam sp_inst_14.INIT_RAM_0A = 256'h1000000400500000000001001100000100040000040040000001100100000100;
defparam sp_inst_14.INIT_RAM_0B = 256'h0040014040400004014050001004100100140400040000000001000000000010;
defparam sp_inst_14.INIT_RAM_0C = 256'h1004000040141010000000000001005410140000000000004015014000000000;
defparam sp_inst_14.INIT_RAM_0D = 256'h0000001001000104410010010040040100400410000400100001010140110000;
defparam sp_inst_14.INIT_RAM_0E = 256'h0110004001000400100040010004001000400100040100040400400004000400;
defparam sp_inst_14.INIT_RAM_0F = 256'h0000000000000000004004000411044500040000000001140010000000000401;
defparam sp_inst_14.INIT_RAM_10 = 256'h0000010000010000000000004004000004000100010000400010004000004000;
defparam sp_inst_14.INIT_RAM_11 = 256'h4004010010040100104000100040000404050044000040040004110400400100;
defparam sp_inst_14.INIT_RAM_12 = 256'h0004001000400100040010004001000400100400101001000010001000000000;
defparam sp_inst_14.INIT_RAM_13 = 256'h0100100010001011011044111400100000000004500040000000001004044001;
defparam sp_inst_14.INIT_RAM_14 = 256'h0000040100004014041410000400000040040004004000400004000100004000;
defparam sp_inst_14.INIT_RAM_15 = 256'h0041000100000000000000000000000000000400000100044010010040000401;
defparam sp_inst_14.INIT_RAM_16 = 256'h4000040000101000100451000040000000010000001000040001000100000410;
defparam sp_inst_14.INIT_RAM_17 = 256'h0000000400010000001000000400001004000040000101000100000040000100;
defparam sp_inst_14.INIT_RAM_18 = 256'h0000000004000000100000000100000100000001000100000000000010000400;
defparam sp_inst_14.INIT_RAM_19 = 256'h1000001000100040000000000100400010000000000000000400000000400001;
defparam sp_inst_14.INIT_RAM_1A = 256'h0100000400004040040004000010000500011000001000000040001000004000;
defparam sp_inst_14.INIT_RAM_1B = 256'h0040104011004000000000401104100440410044010001040110040000000000;
defparam sp_inst_14.INIT_RAM_1C = 256'h0000000010001004000001000400001010004000004000110104011004100440;
defparam sp_inst_14.INIT_RAM_1D = 256'h0000010001001000000000000000000000000100000000000000001000000000;
defparam sp_inst_14.INIT_RAM_1E = 256'h0100000000000000040000000000000010000010000010000000004000000001;
defparam sp_inst_14.INIT_RAM_1F = 256'h4004000110400000101001004410050000000100000100000000040100100100;
defparam sp_inst_14.INIT_RAM_20 = 256'h4004000100100100000000000000040000000000010000000000000040100000;
defparam sp_inst_14.INIT_RAM_21 = 256'h1000001000000000004010000000400000000001001040000400000001000000;
defparam sp_inst_14.INIT_RAM_22 = 256'h0000014000000000004400010051000000400000110504000100001001000000;
defparam sp_inst_14.INIT_RAM_23 = 256'h1040004040010001010004000404001000101040004000401000505044000044;
defparam sp_inst_14.INIT_RAM_24 = 256'h4410400010010010000400104040104040110410000400050400040410001014;
defparam sp_inst_14.INIT_RAM_25 = 256'h0400004004011040001000004004011040001001001000010000410100410100;
defparam sp_inst_14.INIT_RAM_26 = 256'h0100004100010105410001041000104100010414104000404010100401004000;
defparam sp_inst_14.INIT_RAM_27 = 256'h0404410004004004000000000441000400100100040041010440040110400010;
defparam sp_inst_14.INIT_RAM_28 = 256'h0040110040104400154100001000500401044104400000100100100404410010;
defparam sp_inst_14.INIT_RAM_29 = 256'h0004040040040110444100004004410550000100054100001000441400100414;
defparam sp_inst_14.INIT_RAM_2A = 256'h4000040041404414044140440400401104000100100040110504000040040000;
defparam sp_inst_14.INIT_RAM_2B = 256'h4000400004410440011041041100000000400004001104100004005040110441;
defparam sp_inst_14.INIT_RAM_2C = 256'h0000044101104104104411001000100010001000100010004000400040004000;
defparam sp_inst_14.INIT_RAM_2D = 256'h1044110010001000100010001000100040004000400040000441044001400000;
defparam sp_inst_14.INIT_RAM_2E = 256'h0004001001000000001010410001104000000100440010000000044101104104;
defparam sp_inst_14.INIT_RAM_2F = 256'h1104000100100401000000040010004010441000040040400010010401105040;
defparam sp_inst_14.INIT_RAM_30 = 256'h0400000000000040110410404001104104040040000100100040000000040040;
defparam sp_inst_14.INIT_RAM_31 = 256'h0000000004000044100000004000000400050441000041004410000400000010;
defparam sp_inst_14.INIT_RAM_32 = 256'h0100110510510100441000040040040010400104100000010000001001040001;
defparam sp_inst_14.INIT_RAM_33 = 256'h1010040110400010010400400104000000004010100401104000100100040000;
defparam sp_inst_14.INIT_RAM_34 = 256'h4011000400000010010044040110400010010400410014000000100000110000;
defparam sp_inst_14.INIT_RAM_35 = 256'h0000400410010400500000004000004400004041040041000400000000401010;
defparam sp_inst_14.INIT_RAM_36 = 256'h0110010000001000044000000044000044000100000400400100100000010401;
defparam sp_inst_14.INIT_RAM_37 = 256'h1000010040400004010100001004040000401010000100404000040101000010;
defparam sp_inst_14.INIT_RAM_38 = 256'h0004010100001004040000401010000100404000040101000010040400004010;
defparam sp_inst_14.INIT_RAM_39 = 256'h1004040000401010000100404000040101000010040400004010100001004040;
defparam sp_inst_14.INIT_RAM_3A = 256'h1010000100404000040101000010040400004010100001004040000401010000;
defparam sp_inst_14.INIT_RAM_3B = 256'h4000000100000010040400004010100001004040000401010000100404000040;
defparam sp_inst_14.INIT_RAM_3C = 256'h0404100040000000001000000040100000000000000100400000100400400100;
defparam sp_inst_14.INIT_RAM_3D = 256'h0000000000000000050140141004000001001000400041044440000100100001;
defparam sp_inst_14.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3F = 256'h5154455010154040110104445114000001144405140511400115151550054000;

SP sp_inst_15 (
    .DO({sp_inst_15_dout_w[15:0],sp_inst_15_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_15.READ_MODE = 1'b0;
defparam sp_inst_15.WRITE_MODE = 2'b01;
defparam sp_inst_15.BIT_WIDTH = 16;
defparam sp_inst_15.BLK_SEL = 3'b001;
defparam sp_inst_15.RESET_MODE = "SYNC";
defparam sp_inst_15.INIT_RAM_00 = 256'h613C6D5B346D006562206572612069642D2D3E6561763E72613C6D5B316D7473;
defparam sp_inst_15.INIT_RAM_01 = 256'h745B00686F7400002D2D765B0076006477206572612069642D2D3E6561763E72;
defparam sp_inst_15.INIT_RAM_02 = 256'h00796564005D6574656D2065635B656D616C000073657265745B000070686863;
defparam sp_inst_15.INIT_RAM_03 = 256'h64775D747420725B00006164005D65747565775B70756177000073657961645B;
defparam sp_inst_15.INIT_RAM_04 = 256'h00003269656C736520632D2D005D6C6165722070695B000032695D747420775B;
defparam sp_inst_15.INIT_RAM_05 = 256'h2072695B00003269746920632D2D3E6164773E7261673C20646469682077695B;
defparam sp_inst_15.INIT_RAM_06 = 256'h625B7465616200632D2D005D615B6461646120632D2D3E7261673C2064646968;
defparam sp_inst_15.INIT_RAM_07 = 256'h5D79635B006D695F6F63005D616C6E696873665F735B00006F6300006E3C6564;
defparam sp_inst_15.INIT_RAM_08 = 256'h736170735D74695F735B7469707374692074755B0074697500003C2064742D2D;
defparam sp_inst_15.INIT_RAM_09 = 256'h735B687366735D64725F735B000070736574775F735B000070736573655F735B;
defparam sp_inst_15.INIT_RAM_0A = 256'h7F807F78444C7F705D4C4E5B0000554E00745D69655B0000695F70676873665F;
defparam sp_inst_15.INIT_RAM_0B = 256'h801C80084ADC80047FF87FE444747FDC7FC87FB449BC7FB07F9C7F8848A87F84;
defparam sp_inst_15.INIT_RAM_0C = 256'h806C808C53408084806C807C508C8074806C80684E0C8064804C80384B6C8034;
defparam sp_inst_15.INIT_RAM_0D = 256'h806C80F056C880E8806C80D855D880D0806C80C054D480B8806C80A45440809C;
defparam sp_inst_15.INIT_RAM_0E = 256'h819481785FC48170816481405EB88138812881145E6C810C806C81005DE880FC;
defparam sp_inst_15.INIT_RAM_0F = 256'h820081F86CD481EC806C81D463B881CC806C81BC624881B481AC81A460A481A0;
defparam sp_inst_15.INIT_RAM_10 = 256'h806C8254665C824C806C824068FC8238806C822C65F48224806C821865488210;
defparam sp_inst_15.INIT_RAM_11 = 256'h806C82946CA8829C806C82946C748288806C827C698C8274806C8268678C8260;
defparam sp_inst_15.INIT_RAM_12 = 256'h4F52090A73252509090A0D0A3A64200900003A73616D630A82A082A8488882A0;
defparam sp_inst_15.INIT_RAM_13 = 256'h000042410A0D240A0D0A6D63207068206761200A000A21646D6D206566657520;
defparam sp_inst_15.INIT_RAM_14 = 256'h3E6D3C2072643C2064206761200A0A0D203D756E0A0D203D656C0D733D207473;
defparam sp_inst_15.INIT_RAM_15 = 256'h00093830300A0D0A756E3E72613C64206761200A20782520093A3025200A0000;
defparam sp_inst_15.INIT_RAM_16 = 256'h61763E72613C6D206761200A00003E6561763E72613C6D206761200A20782520;
defparam sp_inst_15.INIT_RAM_17 = 256'h76206761200A0A2E7265756E61676C690A2E7265756E656861676C6900003E65;
defparam sp_inst_15.INIT_RAM_18 = 256'h652065746120642050560A20747273206574612064205056000D6D75203E6461;
defparam sp_inst_15.INIT_RAM_19 = 256'h6C6F535478383020202063735354783830202020727453540A3A736E540A000A;
defparam sp_inst_15.INIT_RAM_1A = 256'h302020787830205D255B000065524320202072746E6820202020783830206D69;
defparam sp_inst_15.INIT_RAM_1B = 256'h20392020202030203630203520202020302032302031202020202020200A7838;
defparam sp_inst_15.INIT_RAM_1C = 256'h6E773C206E696375200A00006E696176630A000025206C616162000031203031;
defparam sp_inst_15.INIT_RAM_1D = 256'h6F446375200A00006F64000063536375200A0000637300006E496375200A3E68;
defparam sp_inst_15.INIT_RAM_1E = 256'h002E6F506375200A00006F700000656E68633E686E773C206F646375200A6854;
defparam sp_inst_15.INIT_RAM_1F = 256'h202020200920745F6F64746920686F746567550A2E7272457570200A00006873;
defparam sp_inst_15.INIT_RAM_20 = 256'h200A206E7320756F2020202020202020203E6E6E633C6874776F206E6420756F;
defparam sp_inst_15.INIT_RAM_21 = 256'h00002E2E72612072697465700A0D6F686863742020200A096C6C20686F742020;
defparam sp_inst_15.INIT_RAM_22 = 256'h726120726974726F0A0D3E633C206D5F6174203E646F65707465203A61730A0D;
defparam sp_inst_15.INIT_RAM_23 = 256'h73753A656D3C616C203A61730A0D636520726974203A61730A0D642567722E2E;
defparam sp_inst_15.INIT_RAM_24 = 256'h2E74747355206157656D0A0D00730A0D736D0A0D73750A0D3E6C3C203A336D3A;
defparam sp_inst_15.INIT_RAM_25 = 256'h0A0D65626E20206561726E6F0A0D3E633C20656B203A61730A0D000A3A63612E;
defparam sp_inst_15.INIT_RAM_26 = 256'h732020736D6D68202D6D79792D2061640000202E6974616C6964742061640A0D;
defparam sp_inst_15.INIT_RAM_27 = 256'h7A482D20616400002E742074206F73736D3A20646D6D2D20616400002E657420;
defparam sp_inst_15.INIT_RAM_28 = 256'h65746172206B686300002E6563737020732020726574206E7963716520746E69;
defparam sp_inst_15.INIT_RAM_29 = 256'h6F662D2061640D7A3836332020656C636220756F0A0D006D6170696C6E69000A;
defparam sp_inst_15.INIT_RAM_2A = 256'h8AAC662D692D732D682D64323A64253A3025002030253230643230320D657375;
defparam sp_inst_15.INIT_RAM_2B = 256'h63652067203A61730A0D0000253A72612E2E6174747320670A0D8AB88AB48AB0;
defparam sp_inst_15.INIT_RAM_2C = 256'h303D646178253D6164773E6164773E7261673C2064646968207769206761200A;
defparam sp_inst_15.INIT_RAM_2D = 256'h0A0D000A3230302061640A0D000A64646572726470693C7269206761200A0078;
defparam sp_inst_15.INIT_RAM_2E = 256'h2C5052562820495F4129202C5F4329303A6C0A0D003E6D69203E643C6C652043;
defparam sp_inst_15.INIT_RAM_2F = 256'h203A3A760A0D636D6164282065723628293128563129202C4F52342856302933;
defparam sp_inst_15.INIT_RAM_30 = 256'h2C305047202C5F4320306E3C656462206761200A00647461636C0A0D6420202C;
defparam sp_inst_15.INIT_RAM_31 = 256'h2F31746975206761200A726F65206F63002E0072656D61706E6F0A0D314F4720;
defparam sp_inst_15.INIT_RAM_32 = 256'h202E0A7474737469200A00003E72613C746973206761200A0D78303D0A0D0A20;
defparam sp_inst_15.INIT_RAM_33 = 256'h6174722072726B63630A000A61746461200A203E6461646173206761200A000A;
defparam sp_inst_15.INIT_RAM_34 = 256'h617272700A7474737361200A00003E72613C736173206761200A782564642078;
defparam sp_inst_15.INIT_RAM_35 = 256'h0A0D000A6F6463650A0D000A6174747563650A0D656E206D676F0A0D0A747473;
defparam sp_inst_15.INIT_RAM_36 = 256'h73256E756425656E20200A0D0000252C2C78726F65206F630A0D61746D617970;
defparam sp_inst_15.INIT_RAM_37 = 256'h4B3A49686F742D0A0D0A2E2E2E2E2E2E544E54462E2E2E2E2E2E2E0A00003E20;
defparam sp_inst_15.INIT_RAM_38 = 256'h2E2E2E0A0D0A2E2E2E2E2E2E4C495F542E2E2E2E2E2E2E0A000A7830656E6843;
defparam sp_inst_15.INIT_RAM_39 = 256'h2E7472726E696165207269546C6168706550000D2E2E2E2E2E2E2E432E2E2E2E;
defparam sp_inst_15.INIT_RAM_3A = 256'h6E586E0C000A747072656920656C726554206F43000025787663203161750000;
defparam sp_inst_15.INIT_RAM_3B = 256'h731872CC7280723471E8719C7150710470B8706C70206FD46F886F3C6EF06EA4;
defparam sp_inst_15.INIT_RAM_3C = 256'h79DC7A2C774076F476A8765C761075C47578752C74E07494744873FC73B07364;
defparam sp_inst_15.INIT_RAM_3D = 256'h786579F87A2C7A2C7A2C7A2C7A2C7A2C7A2C7A2C7A2C7A2C7A2C7A2C7A2C7A2C;
defparam sp_inst_15.INIT_RAM_3E = 256'h61687269616F675F7865656C61687269616F675F7865656C61687269616F675F;
defparam sp_inst_15.INIT_RAM_3F = 256'h616F675F7865656C61687269616F675F7865656C61687269616F675F7865656C;

SP sp_inst_16 (
    .DO({sp_inst_16_dout_w[15:0],sp_inst_16_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_16.READ_MODE = 1'b0;
defparam sp_inst_16.WRITE_MODE = 2'b01;
defparam sp_inst_16.BIT_WIDTH = 16;
defparam sp_inst_16.BLK_SEL = 3'b001;
defparam sp_inst_16.RESET_MODE = "SYNC";
defparam sp_inst_16.INIT_RAM_00 = 256'h646420340000000074797373646479666F6D005D756C3C206464203100000000;
defparam sp_inst_16.INIT_RAM_01 = 256'h756F0000637500003176005D00000000726F7373646479666F6D005D756C3C20;
defparam sp_inst_16.INIT_RAM_02 = 256'h0000616C0000747320726974726F0072697400005D7474206D6900007465005D;
defparam sp_inst_16.INIT_RAM_03 = 256'h0067000073656374000065740000747320706B610000656B00005D7474206C65;
defparam sp_inst_16.INIT_RAM_04 = 256'h00007763000061637270326900003E656373703C633200007063000073656764;
defparam sp_inst_16.INIT_RAM_05 = 256'h633C633200007263006572773269005D74613C20646465723E726170633C6332;
defparam sp_inst_16.INIT_RAM_06 = 256'h74610000647400006461000063640063000065723269005D646465723E726170;
defparam sp_inst_16.INIT_RAM_07 = 256'h0000706F00006172797000006873665F3E3D616C69700000797000005D3E2074;
defparam sp_inst_16.INIT_RAM_08 = 256'h006572650000696E697000006E69005D6E6972610000696E00003E6E74656162;
defparam sp_inst_16.INIT_RAM_09 = 256'h69700000616C00006165697000006472005D6972697000007277005D61726970;
defparam sp_inst_16.INIT_RAM_0A = 256'h1C001C001C001C0000004C5500004C4C0000000074780000746E6F69005D616C;
defparam sp_inst_16.INIT_RAM_0B = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_0C = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_0D = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_0E = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_0F = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_10 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_11 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_12 = 256'h3A525245000A0973732500007325322500000A0A646E6D6F1C001C001C001C00;
defparam sp_inst_16.INIT_RAM_13 = 256'h000044430000002000003E643C206C653A657375000021216E616F636E69646E;
defparam sp_inst_16.INIT_RAM_14 = 256'h0D0A756E203E646120313A65737500006425206D00006425206E000A25203072;
defparam sp_inst_16.INIT_RAM_15 = 256'h00003A78257800003E6D3C20646420343A657375000032300000783878300000;
defparam sp_inst_16.INIT_RAM_16 = 256'h756C3C20646420343A65737500000D0A756C3C20646420313A65737500003830;
defparam sp_inst_16.INIT_RAM_17 = 256'h3C203A65737500002E2E626D206C656C00002E2E626D2078206C656C00000D0A;
defparam sp_inst_16.INIT_RAM_18 = 256'h646E74732064616D4D5700006465617474732064616D4D5700000A3E6E3C7264;
defparam sp_inst_16.INIT_RAM_19 = 256'h546C505F000A25783D2068544F5F000A25783D20206C435F0000726F65730000;
defparam sp_inst_16.INIT_RAM_1A = 256'h257820203825203D643200000A73746E20202020744143202020000A25783D20;
defparam sp_inst_16.INIT_RAM_1B = 256'h202030203830203720202020302034302033202020203020303020202020000A;
defparam sp_inst_16.INIT_RAM_1C = 256'h745F6F64746920686F7400007469006C746E000064340000767300000A312020;
defparam sp_inst_16.INIT_RAM_1D = 256'h6E7720686F5400006E7700006E6120686F5400006E610000746920686F54002E;
defparam sp_inst_16.INIT_RAM_1E = 256'h00006C6C20686F5400006C6C00003E6C6E613C20745F6F646E7720686F740000;
defparam sp_inst_16.INIT_RAM_1F = 256'h742020200A093E686E773C206E696375203A617300006F7220746E490000776F;
defparam sp_inst_16.INIT_RAM_20 = 256'h2020090961636863742020200A20202020096C656168203E5F6E643C776F6863;
defparam sp_inst_16.INIT_RAM_21 = 256'h00000A2E2E747473656D2074682000777320756F2020202009206F7063752020;
defparam sp_inst_16.INIT_RAM_22 = 256'h2E747473656D20656320000065733E737472733C636969723C20706865675520;
defparam sp_inst_16.INIT_RAM_23 = 256'h322C3A31646F2079656465675520003E733C656D616C65675520000A3A63612E;
defparam sp_inst_16.INIT_RAM_24 = 256'h2E2E72612070656B20726954000064250000642500006425000061763E732C73;
defparam sp_inst_16.INIT_RAM_25 = 256'h000021726D75666F676E20677277000065737075617765675520000064256772;
defparam sp_inst_16.INIT_RAM_26 = 256'h74656F74733A3A6864646D2D2073657400000A0D656D20797073206F65740000;
defparam sp_inst_16.INIT_RAM_27 = 256'h3A202066657400000A0D6E69657374203A6D6868642D2069657400000A0D6D69;
defparam sp_inst_16.INIT_RAM_28 = 256'h0D72656D6170636500000A0D6C61657274656F7465676E6969206E6572667570;
defparam sp_inst_16.INIT_RAM_29 = 256'h207220686574000A482037326F74736F2065646C687300006172206461760000;
defparam sp_inst_16.INIT_RAM_2A = 256'h1C0000000000000000000000302532306432000064322D64252D3025000A6761;
defparam sp_inst_16.INIT_RAM_2B = 256'h003E733C64776567552000000A6463672E2E74727320657464771C001C001C00;
defparam sp_inst_16.INIT_RAM_2C = 256'h25787264000078307461000A74613C20646465723E726170633C63323A657375;
defparam sp_inst_16.INIT_RAM_2D = 256'h444100000D7825786174722000003E7261673C3E6461686363323A6573750000;
defparam sp_inst_16.INIT_RAM_2E = 256'h2820414329322C3143443128304944412820657300007365743C7669203E733C;
defparam sp_inst_16.INIT_RAM_2F = 256'h3264302069640000616329372C667629202C7276302E352854555629202C2E31;
defparam sp_inst_16.INIT_RAM_30 = 256'h32204F49203130494441203E207474613A657375000025656C75616300343A31;
defparam sp_inst_16.INIT_RAM_31 = 256'h3E323C206E693A657375000A72727970000000006574617220677277000A4950;
defparam sp_inst_16.INIT_RAM_32 = 256'h0000000072612065727700000A206464206572773A657375000A257864690000;
defparam sp_inst_16.INIT_RAM_33 = 256'h253D6164726F652065680000747273206572000A72643C2065723A6573750000;
defparam sp_inst_16.INIT_RAM_34 = 256'h206D676F000072612065726500000A206464206572653A657375000A3D726169;
defparam sp_inst_16.INIT_RAM_35 = 256'h6F630000656E206B68630000747273206F6B6863000A6F646172727000007261;
defparam sp_inst_16.INIT_RAM_36 = 256'h20203A636620203A696C3C2000000A7878252520727279700000747273207269;
defparam sp_inst_16.INIT_RAM_37 = 256'h7965746E63752D2D00002E2E2E2E2E2E2E2E495F4F532E2E2E2E2E2E00000A0D;
defparam sp_inst_16.INIT_RAM_38 = 256'h2E2E2E2E00002E2E2E2E2E2E2E2E414641422E2E2E2E2E2E000078253A6C6E61;
defparam sp_inst_16.INIT_RAM_39 = 256'h0A2E7075657420726C63656D20737265697200000A2E2E2E2E2E2E2E44412E2E;
defparam sp_inst_16.INIT_RAM_3A = 256'h1C001C0000002E2E7572746E726163206D69657200000A78303A657274720000;
defparam sp_inst_16.INIT_RAM_3B = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_3C = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_3D = 256'h69741C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_16.INIT_RAM_3E = 256'h646E5F715F32697069740072646E5F715F31697069740072646E5F715F306970;
defparam sp_inst_16.INIT_RAM_3F = 256'h5F35697069740072646E5F715F34697069740072646E5F715F33697069740072;

SP sp_inst_17 (
    .DO(sp_inst_17_dout[31:0]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[8:0],gw_gnd,gw_vcc,gw_vcc,gw_vcc,gw_vcc}),
    .DI(din[31:0])
);

defparam sp_inst_17.READ_MODE = 1'b0;
defparam sp_inst_17.WRITE_MODE = 2'b01;
defparam sp_inst_17.BIT_WIDTH = 32;
defparam sp_inst_17.BLK_SEL = 3'b001;
defparam sp_inst_17.RESET_MODE = "SYNC";
defparam sp_inst_17.INIT_RAM_00 = 256'h646E61685F7172695F36616F6970675F697478650072656C646E61685F717269;
defparam sp_inst_17.INIT_RAM_01 = 256'h697478650072656C646E61685F7172695F37616F6970675F697478650072656C;
defparam sp_inst_17.INIT_RAM_02 = 256'h5F31626F6970675F697478650072656C646E61685F7172695F30626F6970675F;
defparam sp_inst_17.INIT_RAM_03 = 256'h646E61685F7172695F32626F6970675F697478650072656C646E61685F717269;
defparam sp_inst_17.INIT_RAM_04 = 256'h697478650072656C646E61685F7172695F33626F6970675F697478650072656C;
defparam sp_inst_17.INIT_RAM_05 = 256'h5F35626F6970675F697478650072656C646E61685F7172695F34626F6970675F;
defparam sp_inst_17.INIT_RAM_06 = 256'h646E61685F7172695F36626F6970675F697478650072656C646E61685F717269;
defparam sp_inst_17.INIT_RAM_07 = 256'h697478650072656C646E61685F7172695F37626F6970675F697478650072656C;
defparam sp_inst_17.INIT_RAM_08 = 256'h5F31636F6970675F697478650072656C646E61685F7172695F30636F6970675F;
defparam sp_inst_17.INIT_RAM_09 = 256'h646E61685F7172695F32636F6970675F697478650072656C646E61685F717269;
defparam sp_inst_17.INIT_RAM_0A = 256'h697478650072656C646E61685F7172695F33636F6970675F697478650072656C;
defparam sp_inst_17.INIT_RAM_0B = 256'h5F35636F6970675F697478650072656C646E61685F7172695F34636F6970675F;
defparam sp_inst_17.INIT_RAM_0C = 256'h646E61685F7172695F36636F6970675F697478650072656C646E61685F717269;
defparam sp_inst_17.INIT_RAM_0D = 256'h697478650072656C646E61685F7172695F37636F6970675F697478650072656C;
defparam sp_inst_17.INIT_RAM_0E = 256'h5F31646F6970675F697478650072656C646E61685F7172695F30646F6970675F;
defparam sp_inst_17.INIT_RAM_0F = 256'h646E61685F7172695F32646F6970675F697478650072656C646E61685F717269;
defparam sp_inst_17.INIT_RAM_10 = 256'h697478650072656C646E61685F7172695F33646F6970675F697478650072656C;
defparam sp_inst_17.INIT_RAM_11 = 256'h5F35646F6970675F697478650072656C646E61685F7172695F34646F6970675F;
defparam sp_inst_17.INIT_RAM_12 = 256'h646E61685F7172695F36646F6970675F697478650072656C646E61685F717269;
defparam sp_inst_17.INIT_RAM_13 = 256'h5F7478650072656C646E61685F7172695F37646F6970675F697478650072656C;
defparam sp_inst_17.INIT_RAM_14 = 256'h0000000000000000000000001C007B601C007B69000000000072656C646E6168;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[10]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(sp_inst_15_dout[0]),
  .I1(sp_inst_17_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(spx9_inst_0_dout[0]),
  .I1(spx9_inst_1_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(spx9_inst_2_dout[0]),
  .I1(spx9_inst_3_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(mux_o_11),
  .I1(mux_o_12),
  .S0(dff_q_1)
);
MUX2 mux_inst_16 (
  .O(dout[0]),
  .I0(mux_o_14),
  .I1(mux_o_10),
  .S0(dff_q_0)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(sp_inst_15_dout[1]),
  .I1(sp_inst_17_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(spx9_inst_0_dout[1]),
  .I1(spx9_inst_1_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(spx9_inst_2_dout[1]),
  .I1(spx9_inst_3_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_1)
);
MUX2 mux_inst_33 (
  .O(dout[1]),
  .I0(mux_o_31),
  .I1(mux_o_27),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(sp_inst_15_dout[2]),
  .I1(sp_inst_17_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(spx9_inst_0_dout[2]),
  .I1(spx9_inst_1_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(spx9_inst_2_dout[2]),
  .I1(spx9_inst_3_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_1)
);
MUX2 mux_inst_50 (
  .O(dout[2]),
  .I0(mux_o_48),
  .I1(mux_o_44),
  .S0(dff_q_0)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(sp_inst_15_dout[3]),
  .I1(sp_inst_17_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(spx9_inst_0_dout[3]),
  .I1(spx9_inst_1_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(spx9_inst_2_dout[3]),
  .I1(spx9_inst_3_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(dff_q_1)
);
MUX2 mux_inst_67 (
  .O(dout[3]),
  .I0(mux_o_65),
  .I1(mux_o_61),
  .S0(dff_q_0)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(sp_inst_15_dout[4]),
  .I1(sp_inst_17_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(spx9_inst_0_dout[4]),
  .I1(spx9_inst_1_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(spx9_inst_2_dout[4]),
  .I1(spx9_inst_3_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_1)
);
MUX2 mux_inst_84 (
  .O(dout[4]),
  .I0(mux_o_82),
  .I1(mux_o_78),
  .S0(dff_q_0)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(sp_inst_15_dout[5]),
  .I1(sp_inst_17_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(spx9_inst_0_dout[5]),
  .I1(spx9_inst_1_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(spx9_inst_2_dout[5]),
  .I1(spx9_inst_3_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(dff_q_1)
);
MUX2 mux_inst_101 (
  .O(dout[5]),
  .I0(mux_o_99),
  .I1(mux_o_95),
  .S0(dff_q_0)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(sp_inst_15_dout[6]),
  .I1(sp_inst_17_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(spx9_inst_0_dout[6]),
  .I1(spx9_inst_1_dout[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(spx9_inst_2_dout[6]),
  .I1(spx9_inst_3_dout[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(dff_q_1)
);
MUX2 mux_inst_118 (
  .O(dout[6]),
  .I0(mux_o_116),
  .I1(mux_o_112),
  .S0(dff_q_0)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(sp_inst_15_dout[7]),
  .I1(sp_inst_17_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(spx9_inst_0_dout[7]),
  .I1(spx9_inst_1_dout[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(spx9_inst_2_dout[7]),
  .I1(spx9_inst_3_dout[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_1)
);
MUX2 mux_inst_135 (
  .O(dout[7]),
  .I0(mux_o_133),
  .I1(mux_o_129),
  .S0(dff_q_0)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(sp_inst_15_dout[8]),
  .I1(sp_inst_17_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(spx9_inst_0_dout[8]),
  .I1(spx9_inst_1_dout[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(spx9_inst_2_dout[8]),
  .I1(spx9_inst_3_dout[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(dff_q_1)
);
MUX2 mux_inst_152 (
  .O(dout[8]),
  .I0(mux_o_150),
  .I1(mux_o_146),
  .S0(dff_q_0)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(sp_inst_15_dout[9]),
  .I1(sp_inst_17_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(spx9_inst_4_dout[9]),
  .I1(spx9_inst_5_dout[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(spx9_inst_6_dout[9]),
  .I1(spx9_inst_7_dout[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(mux_o_164),
  .I1(mux_o_165),
  .S0(dff_q_1)
);
MUX2 mux_inst_169 (
  .O(dout[9]),
  .I0(mux_o_167),
  .I1(mux_o_163),
  .S0(dff_q_0)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(sp_inst_15_dout[10]),
  .I1(sp_inst_17_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(spx9_inst_4_dout[10]),
  .I1(spx9_inst_5_dout[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(spx9_inst_6_dout[10]),
  .I1(spx9_inst_7_dout[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_1)
);
MUX2 mux_inst_186 (
  .O(dout[10]),
  .I0(mux_o_184),
  .I1(mux_o_180),
  .S0(dff_q_0)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(sp_inst_15_dout[11]),
  .I1(sp_inst_17_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(spx9_inst_4_dout[11]),
  .I1(spx9_inst_5_dout[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(spx9_inst_6_dout[11]),
  .I1(spx9_inst_7_dout[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_1)
);
MUX2 mux_inst_203 (
  .O(dout[11]),
  .I0(mux_o_201),
  .I1(mux_o_197),
  .S0(dff_q_0)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(sp_inst_15_dout[12]),
  .I1(sp_inst_17_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(spx9_inst_4_dout[12]),
  .I1(spx9_inst_5_dout[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(spx9_inst_6_dout[12]),
  .I1(spx9_inst_7_dout[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_215),
  .I1(mux_o_216),
  .S0(dff_q_1)
);
MUX2 mux_inst_220 (
  .O(dout[12]),
  .I0(mux_o_218),
  .I1(mux_o_214),
  .S0(dff_q_0)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(sp_inst_15_dout[13]),
  .I1(sp_inst_17_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(spx9_inst_4_dout[13]),
  .I1(spx9_inst_5_dout[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(spx9_inst_6_dout[13]),
  .I1(spx9_inst_7_dout[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_232),
  .I1(mux_o_233),
  .S0(dff_q_1)
);
MUX2 mux_inst_237 (
  .O(dout[13]),
  .I0(mux_o_235),
  .I1(mux_o_231),
  .S0(dff_q_0)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(sp_inst_15_dout[14]),
  .I1(sp_inst_17_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(spx9_inst_4_dout[14]),
  .I1(spx9_inst_5_dout[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(spx9_inst_6_dout[14]),
  .I1(spx9_inst_7_dout[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(mux_o_249),
  .I1(mux_o_250),
  .S0(dff_q_1)
);
MUX2 mux_inst_254 (
  .O(dout[14]),
  .I0(mux_o_252),
  .I1(mux_o_248),
  .S0(dff_q_0)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(sp_inst_15_dout[15]),
  .I1(sp_inst_17_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(spx9_inst_4_dout[15]),
  .I1(spx9_inst_5_dout[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(spx9_inst_6_dout[15]),
  .I1(spx9_inst_7_dout[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(dff_q_1)
);
MUX2 mux_inst_271 (
  .O(dout[15]),
  .I0(mux_o_269),
  .I1(mux_o_265),
  .S0(dff_q_0)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(sp_inst_16_dout[16]),
  .I1(sp_inst_17_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(spx9_inst_4_dout[16]),
  .I1(spx9_inst_5_dout[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(spx9_inst_6_dout[16]),
  .I1(spx9_inst_7_dout[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(mux_o_283),
  .I1(mux_o_284),
  .S0(dff_q_1)
);
MUX2 mux_inst_288 (
  .O(dout[16]),
  .I0(mux_o_286),
  .I1(mux_o_282),
  .S0(dff_q_0)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(sp_inst_16_dout[17]),
  .I1(sp_inst_17_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(spx9_inst_4_dout[17]),
  .I1(spx9_inst_5_dout[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(spx9_inst_6_dout[17]),
  .I1(spx9_inst_7_dout[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(dff_q_1)
);
MUX2 mux_inst_305 (
  .O(dout[17]),
  .I0(mux_o_303),
  .I1(mux_o_299),
  .S0(dff_q_0)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(sp_inst_16_dout[18]),
  .I1(sp_inst_17_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_315 (
  .O(dout[18]),
  .I0(sp_inst_8_dout[18]),
  .I1(mux_o_310),
  .S0(dff_q_0)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(sp_inst_16_dout[19]),
  .I1(sp_inst_17_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_325 (
  .O(dout[19]),
  .I0(sp_inst_8_dout[19]),
  .I1(mux_o_320),
  .S0(dff_q_0)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(sp_inst_16_dout[20]),
  .I1(sp_inst_17_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_335 (
  .O(dout[20]),
  .I0(sp_inst_9_dout[20]),
  .I1(mux_o_330),
  .S0(dff_q_0)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(sp_inst_16_dout[21]),
  .I1(sp_inst_17_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_345 (
  .O(dout[21]),
  .I0(sp_inst_9_dout[21]),
  .I1(mux_o_340),
  .S0(dff_q_0)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(sp_inst_16_dout[22]),
  .I1(sp_inst_17_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_355 (
  .O(dout[22]),
  .I0(sp_inst_10_dout[22]),
  .I1(mux_o_350),
  .S0(dff_q_0)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(sp_inst_16_dout[23]),
  .I1(sp_inst_17_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_365 (
  .O(dout[23]),
  .I0(sp_inst_10_dout[23]),
  .I1(mux_o_360),
  .S0(dff_q_0)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(sp_inst_16_dout[24]),
  .I1(sp_inst_17_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_375 (
  .O(dout[24]),
  .I0(sp_inst_11_dout[24]),
  .I1(mux_o_370),
  .S0(dff_q_0)
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(sp_inst_16_dout[25]),
  .I1(sp_inst_17_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_385 (
  .O(dout[25]),
  .I0(sp_inst_11_dout[25]),
  .I1(mux_o_380),
  .S0(dff_q_0)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(sp_inst_16_dout[26]),
  .I1(sp_inst_17_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_395 (
  .O(dout[26]),
  .I0(sp_inst_12_dout[26]),
  .I1(mux_o_390),
  .S0(dff_q_0)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(sp_inst_16_dout[27]),
  .I1(sp_inst_17_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_405 (
  .O(dout[27]),
  .I0(sp_inst_12_dout[27]),
  .I1(mux_o_400),
  .S0(dff_q_0)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(sp_inst_16_dout[28]),
  .I1(sp_inst_17_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_415 (
  .O(dout[28]),
  .I0(sp_inst_13_dout[28]),
  .I1(mux_o_410),
  .S0(dff_q_0)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(sp_inst_16_dout[29]),
  .I1(sp_inst_17_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_425 (
  .O(dout[29]),
  .I0(sp_inst_13_dout[29]),
  .I1(mux_o_420),
  .S0(dff_q_0)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(sp_inst_16_dout[30]),
  .I1(sp_inst_17_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_435 (
  .O(dout[30]),
  .I0(sp_inst_14_dout[30]),
  .I1(mux_o_430),
  .S0(dff_q_0)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(sp_inst_16_dout[31]),
  .I1(sp_inst_17_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_445 (
  .O(dout[31]),
  .I0(sp_inst_14_dout[31]),
  .I1(mux_o_440),
  .S0(dff_q_0)
);
endmodule //Gowin_SP_Instr
