//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.01 (64-bit)
//Part Number: GW5AT-LV138PG484AC2/I1
//Device: GW5AT-138
//Device Version: B
//Created Time: Tue Apr  9 23:22:02 2024

module Gowin_SP_Instr (dout, clk, oce, ce, reset, wre, ad, din);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [11:0] ad;
input [31:0] din;

wire [23:0] sp_inst_0_dout_w;
wire [7:0] sp_inst_0_dout;
wire [23:0] sp_inst_1_dout_w;
wire [15:8] sp_inst_1_dout;
wire [15:0] sp_inst_2_dout_w;
wire [15:0] sp_inst_2_dout;
wire [23:0] sp_inst_3_dout_w;
wire [23:16] sp_inst_3_dout;
wire [23:0] sp_inst_4_dout_w;
wire [31:24] sp_inst_4_dout;
wire [15:0] sp_inst_5_dout_w;
wire [31:16] sp_inst_5_dout;
wire dff_q_0;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],sp_inst_0_dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b01;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h8CEC8C8C2C2C0C2C2CAC8C80ACAD0D8C0CCF8EEF2F8C2CAD0F900FF0EF4F000D;
defparam sp_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000200020006323800C2C8C6C2C;
defparam sp_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_20 = 256'hA08DA08DA08DA08DA08D0CA3A1ABAAA9A8A7A6A5A4B4B3B2B1B0AFAEADAC5535;
defparam sp_inst_0.INIT_RAM_21 = 256'hA5A4B4B3B2B1B0AFAEADAC550000A08D000000000000000000000000A08DA08D;
defparam sp_inst_0.INIT_RAM_22 = 256'hC6C5C4767661632063766100000485CCCC8C767661630015A3A1ABAAA9A8A7A6;
defparam sp_inst_0.INIT_RAM_23 = 256'hCCCC07A0CCCECDACCDCECDCC0780AECDCC00C0CCCC00FF04CC0CCC80CC80CCC7;
defparam sp_inst_0.INIT_RAM_24 = 256'h008C8C8CCC8D0CCDCC0C008CACCD8CCC8DCCCD00CCCC8CCEADCECDCC9FCCCC8C;
defparam sp_inst_0.INIT_RAM_25 = 256'hCCFF84CCFF04AC0CCD00C47676616320637661840C0CCCCC8CCCFF848C8C8CCC;
defparam sp_inst_0.INIT_RAM_26 = 256'h00C0CCCCCC8CCCCBCAC9C8C7C6C5C47676616320637661840C9FCCCC8CCCCC8C;
defparam sp_inst_0.INIT_RAM_27 = 256'hCCCC8CCCFF848CCC808CAC8C2C8DAC0D8C8CACCD8CCCCC0CAC0CCDCC8CACCDCC;
defparam sp_inst_0.INIT_RAM_28 = 256'h078CCC00CC8CCCCC8CCCFF84C506078CCC00CC8CCCCC8CCCFF848C8CCC00CC8C;
defparam sp_inst_0.INIT_RAM_29 = 256'hFF84C506078CCC00CC8CCCCC8CCCFF84C506078CCC00CC8CCCCC8CCCFF84C506;
defparam sp_inst_0.INIT_RAM_2A = 256'h00C0CC8CCC00CC8CCCFF0400CC8CCCCC8CCCFF84C506078CCC00CC8CCCCC8CCC;
defparam sp_inst_0.INIT_RAM_2B = 256'hCD00C0FF8D0C8DACCD8CCC8D0C8DACCD8CCCCC8CCCCCAC8C8CCCCE8CCCAD0CCD;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000FF04FF8D0C8DACCD8CCC8D0C8DACCD8CCCCC8CCCCCAC8C8CCCCE8CCCAD0C;
defparam sp_inst_0.INIT_RAM_2D = 256'h8C8CCC00CCACC476766320637661840C9F8CACCDCCCC8CCCFF84CCFF04AC0CCD;
defparam sp_inst_0.INIT_RAM_2E = 256'hCDC5C4767663206376002C0C7676632063760020767663206376008DCDCC9F8C;
defparam sp_inst_0.INIT_RAM_2F = 256'h80CCCC8CCC008DAD0C8ECCCC0E8D0C008DAD0C8E0CCCCC0E8D0C80CCCCCC8D0C;
defparam sp_inst_0.INIT_RAM_30 = 256'hAD0C8D8C0C767663206376008DAD0C8ECCCC0E8D0C008DAD0C8E0CCCCC0E8D0C;
defparam sp_inst_0.INIT_RAM_31 = 256'h206376008DADAD0C767663206376008DCCADCC8DCCC5C4767663206376008DAD;
defparam sp_inst_0.INIT_RAM_32 = 256'h8C8C0C8DCDCD0C8E0CC476766320637684CCC000CC0C80ACCC8D0CC0C4767663;
defparam sp_inst_0.INIT_RAM_33 = 256'h63FF9FCD8DCC0000000000CC8C6C8DAD0C8D0C767663206376008DADAD8C0C8D;
defparam sp_inst_0.INIT_RAM_34 = 256'h63766100FF840C05FF842405C626767661632063766100FF8DAD0C8D0C767661;
defparam sp_inst_0.INIT_RAM_35 = 256'h0C05FF842405C626767661632063766100FF840C05FF842405C6267676616320;
defparam sp_inst_0.INIT_RAM_36 = 256'hC626767661632063766100FF840C05FF842405C626767661632063766100FF84;
defparam sp_inst_0.INIT_RAM_37 = 256'h2063766100FF840C05FF842405C626767661632063766100FF840C05FF842405;
defparam sp_inst_0.INIT_RAM_38 = 256'h840C05FF842405C626767661632063766100FF840C05FF842405C62676766163;
defparam sp_inst_0.INIT_RAM_39 = 256'h05C626767661632063766100FF840C05FF842405C626767661632063766100FF;
defparam sp_inst_0.INIT_RAM_3A = 256'h632063766100FF840C05FF842405C626767661632063766100FF840C05FF8424;
defparam sp_inst_0.INIT_RAM_3B = 256'hFF840C25FF842405C626767661632063766100FF840C05FF842405C626767661;
defparam sp_inst_0.INIT_RAM_3C = 256'h2405C626767661632063766100FF840C45FF842405C626767661632063766100;
defparam sp_inst_0.INIT_RAM_3D = 256'h61632063766100FF840C05FF842405C626767661632063766100FF840C85FF84;
defparam sp_inst_0.INIT_RAM_3E = 256'h00FF840C05FF842405C626767661632063766100FF840C05FF842405C6267676;
defparam sp_inst_0.INIT_RAM_3F = 256'h842405C626767661632063766100FF840C05FF842405C6267676616320637661;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[23:0],sp_inst_1_dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:8]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b01;
defparam sp_inst_1.BIT_WIDTH = 8;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'hFDE311FD0010003000F911011101000100D135010001001102350235E1002000;
defparam sp_inst_1.INIT_RAM_01 = 256'h000000000000000000000000000000000000000000800008F00001204041A044;
defparam sp_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_20 = 256'h2D812D412D212D1165F114425262728292A2B2C2D2728292A2B2C2D2E2F200C4;
defparam sp_inst_1.INIT_RAM_21 = 256'hC2D2728292A2B2C2D2E2F20004A80D0114141C0824F02CBC34383CF82D012D01;
defparam sp_inst_1.INIT_RAM_22 = 256'h526272C0A0B04000806070008CD001BEBE008060708038C4425262728292A2B2;
defparam sp_inst_1.INIT_RAM_23 = 256'hB2920009359252C135C2B25D0009B1925250B292720C87B49230721D72254242;
defparam sp_inst_1.INIT_RAM_24 = 256'h1481C18182192482820008C131C2FDA21DB2A274A23135B531B2B262B192B205;
defparam sp_inst_1.INIT_RAM_25 = 256'h723301BE3F340D28BE3072C0A0B04000C0A0B001008CA2A2FDA29701815D8182;
defparam sp_inst_1.INIT_RAM_26 = 256'h30B2A272729182726252423222123200E0F08000C0A0B00100C5BEBE01727205;
defparam sp_inst_1.INIT_RAM_27 = 256'hB2A211A2DB0101A2010131E10089AD4C6D01313205B29204E5948E8E013132B2;
defparam sp_inst_1.INIT_RAM_28 = 256'h0401A230B205B2A211A2130192280001A268B205B2A211A20F018101A298B205;
defparam sp_inst_1.INIT_RAM_29 = 256'h6B0192080001A2C0B205B2A211A2A30192200001A2F8B205B2A211A2DB019228;
defparam sp_inst_1.INIT_RAM_2A = 256'h3C92B205B238B205B2D39450B205B2A211A2330192400001A288B205B2A211A2;
defparam sp_inst_1.INIT_RAM_2B = 256'h923C92BB95E401313205B2D9C001313205B2B205B292314101313205B2312892;
defparam sp_inst_1.INIT_RAM_2C = 256'h2400B7943F95E401313205B25DC001313205B2B205B292314101313205B23128;
defparam sp_inst_1.INIT_RAM_2D = 256'h8115B200AE00B28070800080E0F00100C5013132B2B205B28F018E9B340D288E;
defparam sp_inst_1.INIT_RAM_2E = 256'h726272C0B0400040300010044030C000403000044030C00080700001AEB2F181;
defparam sp_inst_1.INIT_RAM_2F = 256'h3162B28172681139D60131B20411D69011B9D6013031B20411D63162B272697C;
defparam sp_inst_1.INIT_RAM_30 = 256'h11D48101D44030C000C0B0005139D60131B20451D62851B9D6013031B20451D6;
defparam sp_inst_1.INIT_RAM_31 = 256'h00403000D1A9B4D64030C00080700031B231A231B2A2B2807080004030000181;
defparam sp_inst_1.INIT_RAM_32 = 256'h010DD40135B2DA01DAB280708000C0B001B2B208B20411B17201DAB272C0B040;
defparam sp_inst_1.INIT_RAM_33 = 256'hC0BFE5B2FDB20000000014B2911C0105E001E0807080008070000181050DD481;
defparam sp_inst_1.INIT_RAM_34 = 256'h402030002F81D604DB0000149000402030C00040203000430105E001E0402030;
defparam sp_inst_1.INIT_RAM_35 = 256'hD61043A0003CF000402030C00040203000E381D6088FD00028C000402030C000;
defparam sp_inst_1.INIT_RAM_36 = 256'h5000402030C000402030004B81D620F77000502000402030C000402030009781;
defparam sp_inst_1.INIT_RAM_37 = 256'h0040203000B381D6805F1000788000402030C00040203000FF81D640AB400064;
defparam sp_inst_1.INIT_RAM_38 = 256'h81D600C7B000A4E000402030C000402030006781D60013E0008CB000402030C0;
defparam sp_inst_1.INIT_RAM_39 = 256'hD04000402030C00040203000CF81D6007B8000B81000402030C000402030001B;
defparam sp_inst_1.INIT_RAM_3A = 256'hC000402030003781D600E32000E87000402030C000402030008381D6002F5000;
defparam sp_inst_1.INIT_RAM_3B = 256'h9F81D6004BC00014D000402030C00040203000EB81D60097F00000A000402030;
defparam sp_inst_1.INIT_RAM_3C = 256'h00403000402030C000402030005381D600FF9000280000402030C00040203000;
defparam sp_inst_1.INIT_RAM_3D = 256'h30C00040203000BB81D601673000586000402030C000402030000781D600B360;
defparam sp_inst_1.INIT_RAM_3E = 256'h002381D604CFD0008CC000402030C000402030006F81D6021B00007490004020;
defparam sp_inst_1.INIT_RAM_3F = 256'h7000BC2000402030C00040203000D781D60883A000A4F000402030C000402030;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[15:0],sp_inst_2_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[11],ad[10]}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b01;
defparam sp_inst_2.BIT_WIDTH = 16;
defparam sp_inst_2.BLK_SEL = 3'b010;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'h50C60026407620763061C063002040632076306100008BFF8184D60C100537FF;
defparam sp_inst_2.INIT_RAM_01 = 256'h20763061C063002040632076306100003FFF8184D60C2005EBFF40840024D405;
defparam sp_inst_2.INIT_RAM_02 = 256'h00204063207630610000F3FF8184D60C40059FFF10840024E80580C600264076;
defparam sp_inst_2.INIT_RAM_03 = 256'h30610000A7FF8184D60C800553FFE0840024FC05B0C60026407620763061C063;
defparam sp_inst_2.INIT_RAM_04 = 256'h8184D60C000507FFB08400241405E0C60026407620763061C063002040632076;
defparam sp_inst_2.INIT_RAM_05 = 256'hBBFF808400242C0510C60026407620763061C063002040632076306100005BFF;
defparam sp_inst_2.INIT_RAM_06 = 256'h440540C60026407620763061C063002040632076306100000FFF8184D60C0005;
defparam sp_inst_2.INIT_RAM_07 = 256'h407620763061C06300204063207630610000C3FF8184D60C00056FFF50840024;
defparam sp_inst_2.INIT_RAM_08 = 256'hC0630020406320763061000077FF8184D60C000523FF208400045C0570C60026;
defparam sp_inst_2.INIT_RAM_09 = 256'h2076306100002BFF8184D60C0005D7FFF08400047405A0C60026407620763061;
defparam sp_inst_2.INIT_RAM_0A = 256'hDFFF8184D60C00058BFFC08400048C05D0C60026407620763061C06300204063;
defparam sp_inst_2.INIT_RAM_0B = 256'h00053FFF90840004A80500C60026407620763061C06300204063207630610000;
defparam sp_inst_2.INIT_RAM_0C = 256'h0004C00530C60026407620763061C0630020406320763061000093FF8184D60C;
defparam sp_inst_2.INIT_RAM_0D = 256'h0026407620763061C0630020406320763061000047FF8184D60C0005F3FF6084;
defparam sp_inst_2.INIT_RAM_0E = 256'h7061806300204063207630610000FBFF8184D60C0005A7FF30840004D80560C6;
defparam sp_inst_2.INIT_RAM_0F = 256'hA2CC318C818CD60C4BFFC0840004880550C60026018D000DF18CD60C80766076;
defparam sp_inst_2.INIT_RAM_10 = 256'h2180058CB1ACB2CCA2CD4000B2C00000A2CCB1AC92CCA2CD92CC018C818CD60C;
defparam sp_inst_2.INIT_RAM_11 = 256'h607670610000BD8D7C0CB2CDB2CC058CB2CC0181018C31AC898CB2CC51AD000D;
defparam sp_inst_2.INIT_RAM_12 = 256'h00001FFFB2CC018C118CD60C018D020DF18CD60C807660767061806300208063;
defparam sp_inst_2.INIT_RAM_13 = 256'hD68CBACCFD8C818CC18C018C118CD68C80766076706180630020806360767061;
defparam sp_inst_2.INIT_RAM_14 = 256'h00040185BACC018D3C0D118CD68C018D040DF18CD60CB6CC3D8C818C018C118C;
defparam sp_inst_2.INIT_RAM_15 = 256'h098CD18C018D080DF18CD60C80767076806300208063607670610000F3FF8084;
defparam sp_inst_2.INIT_RAM_16 = 256'hB2CC7D8CCD8C018C118CD60C80766076706180630020806370760000BECC018C;
defparam sp_inst_2.INIT_RAM_17 = 256'h31ACD18C000C898DB2CC718D400CB2CD018DB5CDF00DF18CD60C018E118CD60C;
defparam sp_inst_2.INIT_RAM_18 = 256'hD60C018E118CD60C0BFF008400043C000180118CD60C27FFD08400040180018C;
defparam sp_inst_2.INIT_RAM_19 = 256'h80766076706180630020806360767061000000000800018DB5CDFDADFEED118C;
defparam sp_inst_2.INIT_RAM_1A = 256'h818C058C018C518CFFCC4980008C63FF00045980058C9ECC9ECC018C158CD40C;
defparam sp_inst_2.INIT_RAM_1B = 256'h03FF9580118C9ECC63FF000487FF50040185018CC18CFFCC018DF18CFFCC018D;
defparam sp_inst_2.INIT_RAM_1C = 256'h040C018D340DD10C1DAC340C82CD82CC018CD10C6C00BECC018C118CD10CA2C0;
defparam sp_inst_2.INIT_RAM_1D = 256'hBECC018C118CD10C018D82CDD10C1000018D280DD10CA2C01980A2CC2C00A2CC;
defparam sp_inst_2.INIT_RAM_1E = 256'h70610000018DFC0D0D8CD40C018D200D0D8CD40C1580218C9ECC919F058CBECC;
defparam sp_inst_2.INIT_RAM_1F = 256'h40632076306100003BFF4FFFA08400046BFF407620763061C063002080636076;
defparam sp_inst_2.INIT_RAM_20 = 256'h15F415F415F4156C167016701670167016701670167016701670167015540020;
defparam sp_inst_2.INIT_RAM_21 = 256'h167016701670167016701670167016701670167015F415F415F415F415F415F4;
defparam sp_inst_2.INIT_RAM_22 = 256'h1670167016701670167016701670167016701670167016701670167016701670;
defparam sp_inst_2.INIT_RAM_23 = 256'h140C14E416701670167016701670167016701670167016701670167016701670;
defparam sp_inst_2.INIT_RAM_24 = 256'h13E016701670151C14AC16701670167016701670167016701670167016701474;
defparam sp_inst_2.INIT_RAM_25 = 256'h1D301CE41C981C4C1C001BB41B681B1C1AD01A841A38151C16701670143C1670;
defparam sp_inst_2.INIT_RAM_26 = 256'h21F021A42158210C20C0207420281FDC1F901F441EF81EAC1E601E141DC81D7C;
defparam sp_inst_2.INIT_RAM_27 = 256'h2E2E2E2E2E0A00003E2073256E756425656E20200A0D236C232022D42288223C;
defparam sp_inst_2.INIT_RAM_28 = 256'h2E0A000A7830656E68434B3A49686F742D0A0D0A2E2E2E2E2E2E544E54462E2E;
defparam sp_inst_2.INIT_RAM_29 = 256'h2E2E2E2E2E432E2E2E2E2E2E2E0A0D0A2E2E2E2E2E2E4C495F542E2E2E2E2E2E;
defparam sp_inst_2.INIT_RAM_2A = 256'h265826582658265826082658000A747072656920656C726554206F43000D2E2E;
defparam sp_inst_2.INIT_RAM_2B = 256'h61687269616F675F786526242658265826582658265826582658265826582658;
defparam sp_inst_2.INIT_RAM_2C = 256'h616F675F7865656C61687269616F675F7865656C61687269616F675F7865656C;
defparam sp_inst_2.INIT_RAM_2D = 256'h7865656C61687269616F675F7865656C61687269616F675F7865656C61687269;
defparam sp_inst_2.INIT_RAM_2E = 256'h61687269626F675F7865656C61687269616F675F7865656C61687269616F675F;
defparam sp_inst_2.INIT_RAM_2F = 256'h626F675F7865656C61687269626F675F7865656C61687269626F675F7865656C;
defparam sp_inst_2.INIT_RAM_30 = 256'h7865656C61687269626F675F7865656C61687269626F675F7865656C61687269;
defparam sp_inst_2.INIT_RAM_31 = 256'h61687269636F675F7865656C61687269626F675F7865656C61687269626F675F;
defparam sp_inst_2.INIT_RAM_32 = 256'h636F675F7865656C61687269636F675F7865656C61687269636F675F7865656C;
defparam sp_inst_2.INIT_RAM_33 = 256'h7865656C61687269636F675F7865656C61687269636F675F7865656C61687269;
defparam sp_inst_2.INIT_RAM_34 = 256'h61687269646F675F7865656C61687269636F675F7865656C61687269636F675F;
defparam sp_inst_2.INIT_RAM_35 = 256'h646F675F7865656C61687269646F675F7865656C61687269646F675F7865656C;
defparam sp_inst_2.INIT_RAM_36 = 256'h7865656C61687269646F675F7865656C61687269646F675F7865656C61687269;
defparam sp_inst_2.INIT_RAM_37 = 256'h00000000656C61687865656C61687269646F675F7865656C61687269646F675F;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[23:0],sp_inst_3_dout[23:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[23:16]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b01;
defparam sp_inst_3.BIT_WIDTH = 8;
defparam sp_inst_3.BLK_SEL = 3'b000;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'hBFFF00BF0000150038FF80800080008000FF10800080008080108010B7380015;
defparam sp_inst_3.INIT_RAM_01 = 256'h000000000000000000000000000000000000000000480019BD0000800688EC06;
defparam sp_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_20 = 256'h0040004000400040006E00BEBEBEBEBEBEBEBEBEBEBFBFBFBFBFBFBFBFBF0000;
defparam sp_inst_3.INIT_RAM_21 = 256'hBEBEBFBFBFBFBFBFBFBFBF000015004100170013001400140014001300600042;
defparam sp_inst_3.INIT_RAM_22 = 256'hBEBEBE818181BE0080808040057F153F3F15808080BF4800BEBEBEBEBEBEBEBE;
defparam sp_inst_3.INIT_RAM_23 = 256'hBFBF2A0021BFBE3E10BFBF002A0021BFBE00BFBFBE00FF80BF11BE00BE00BEBE;
defparam sp_inst_3.INIT_RAM_24 = 256'h00678067BF0080BFBF15003E10BFBFBF00BFBF00BF15131312BFBFBEFFBFBF80;
defparam sp_inst_3.INIT_RAM_25 = 256'hBFFE153FFE8000803F00BF808080BF008181811515FFBFBFBFBFFE15678167BF;
defparam sp_inst_3.INIT_RAM_26 = 256'h03BFBFBFBFBF8080808080808080BF818080BE008080801515FF3F3F00BFBF80;
defparam sp_inst_3.INIT_RAM_27 = 256'hBFBF80BFFE1580BF0080109000400281BF0010BF80BFBF8002803F3F0010BFBF;
defparam sp_inst_3.INIT_RAM_28 = 256'h8080BF02BF80BFBF80BFFD15BF801580BF02BF80BFBF80BFFD156780BF02BF80;
defparam sp_inst_3.INIT_RAM_29 = 256'hFC15BF801580BF01BF80BFBF80BFFC15BF801580BF01BF80BFBF80BFFC15BF80;
defparam sp_inst_3.INIT_RAM_2A = 256'h00BFBF80BF01BF80BFFB8001BF80BFBF80BFFC15BF801580BF01BF80BFBF80BF;
defparam sp_inst_3.INIT_RAM_2B = 256'hBF00BFFDFF800010BF80BFFD800010BF80BFBF80BFBF10BF0010BF80BF1C80BF;
defparam sp_inst_3.INIT_RAM_2C = 256'h0040FA80FDFF800010BF80BFFD800010BF80BFBF80BFBF10BF0010BF80BF1C80;
defparam sp_inst_3.INIT_RAM_2D = 256'h6700BF403F15BF8080BF008180801515FC0010BFBFBF80BFFA153FFA8000803F;
defparam sp_inst_3.INIT_RAM_2E = 256'hBFBFBF8080BF0080804001808080BF00808040018080BF00808040003FBFFF40;
defparam sp_inst_3.INIT_RAM_2F = 256'h00BFBFBFBF0081157F1517BF80817F0081147F151417BF80817F00BFBFBF0080;
defparam sp_inst_3.INIT_RAM_30 = 256'h807F67007F8080BF0080804081157F1517BF80817F0081147F151417BF80817F;
defparam sp_inst_3.INIT_RAM_31 = 256'h0080804080964A7F8080BF0080804080BF15BF80BFBFBF8080BF008080400067;
defparam sp_inst_3.INIT_RAM_32 = 256'h00807F8015BF7F807FBF8080BF00808015BFBF00BF800014BF807FBFBF8080BF;
defparam sp_inst_3.INIT_RAM_33 = 256'hBFFFFFBFBFBF4040404000BFBF0080C07F807F8080BF00808040006780807F67;
defparam sp_inst_3.INIT_RAM_34 = 256'h80808040FE807F80F8BE00808200808080BF0080808040FE80C07F807F808080;
defparam sp_inst_3.INIT_RAM_35 = 256'h7F80F8BB00808000808080BF0080808040FD807F80F8BC00808100808080BF00;
defparam sp_inst_3.INIT_RAM_36 = 256'hBF00808080BF0080808040FD807F80F7BA00808000808080BF0080808040FD80;
defparam sp_inst_3.INIT_RAM_37 = 256'h0080808040FC807F80F7B80080BE00808080BF0080808040FC807F80F7B90080;
defparam sp_inst_3.INIT_RAM_38 = 256'h807F82F6B50080BC00808080BF0080808040FC807F81F7B60080BD00808080BF;
defparam sp_inst_3.INIT_RAM_39 = 256'h80BB00808080BF0080808040FB807F84F6B40080BC00808080BF0080808040FC;
defparam sp_inst_3.INIT_RAM_3A = 256'hBF0080808040FB807F90F5B20080BA00808080BF0080808040FB807F88F6B300;
defparam sp_inst_3.INIT_RAM_3B = 256'hFA807F00F5AF0081B800808080BF0080808040FA807FA0F5B00081B900808080;
defparam sp_inst_3.INIT_RAM_3C = 256'h0081B700808080BF0080808040FA807F00F4AE0081B800808080BF0080808040;
defparam sp_inst_3.INIT_RAM_3D = 256'h80BF0080808040F9807F00F4AC0081B600808080BF0080808040FA807F00F4AD;
defparam sp_inst_3.INIT_RAM_3E = 256'h40F9807F00F3A90081B400808080BF0080808040F9807F00F4AB0081B5008080;
defparam sp_inst_3.INIT_RAM_3F = 256'hA70081B300808080BF0080808040F8807F00F3A80081B300808080BF00808080;

SP sp_inst_4 (
    .DO({sp_inst_4_dout_w[23:0],sp_inst_4_dout[31:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:24]})
);

defparam sp_inst_4.READ_MODE = 1'b0;
defparam sp_inst_4.WRITE_MODE = 2'b01;
defparam sp_inst_4.BIT_WIDTH = 8;
defparam sp_inst_4.BLK_SEL = 3'b000;
defparam sp_inst_4.RESET_MODE = "SYNC";
defparam sp_inst_4.INIT_RAM_00 = 256'h0315040314040004145F022958031503155F0003150315022900280003145000;
defparam sp_inst_4.INIT_RAM_01 = 256'h00000000000000000000000000000000000000004C064C540315040304031404;
defparam sp_inst_4.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_20 = 256'h4403440344034403400304292929292929292929292929292929292929291504;
defparam sp_inst_4.INIT_RAM_21 = 256'h2828282828282828282828155054400350545054505450545054505444034403;
defparam sp_inst_4.INIT_RAM_22 = 256'h292929022929024C022828035415002A29000229290206042828282828282828;
defparam sp_inst_4.INIT_RAM_23 = 256'h2829005C0028282900022800005C002828502929285057022900286428402829;
defparam sp_inst_4.INIT_RAM_24 = 256'h5000020028600228290050280002022860282850290000000028282847282902;
defparam sp_inst_4.INIT_RAM_25 = 256'h2857002A57025C02285029022929024C02282800006328290228570000020028;
defparam sp_inst_4.INIT_RAM_26 = 256'h502929282902022929292929292929022929024C02282800004728292A282902;
defparam sp_inst_4.INIT_RAM_27 = 256'h28290228570028284C2800021C00680202280028022829025C0228292A002828;
defparam sp_inst_4.INIT_RAM_28 = 256'h0228285029022829022857002802002828502902282902285700002828502902;
defparam sp_inst_4.INIT_RAM_29 = 256'h5700280200282850290228290228570028020028285029022829022857002802;
defparam sp_inst_4.INIT_RAM_2A = 256'h5029290228502902285702502902282902285700280200282850290228290228;
defparam sp_inst_4.INIT_RAM_2B = 256'h2850295367022800280228670228002802282902282900022800280228000228;
defparam sp_inst_4.INIT_RAM_2C = 256'h5003570253670228002802286702280028022829022829000228002802280002;
defparam sp_inst_4.INIT_RAM_2D = 256'h002A28032900290229024C0228280000472800282829022857002A57025C0228;
defparam sp_inst_4.INIT_RAM_2E = 256'h2829290229024C02280304030229024C022803040229024C022803292A284303;
defparam sp_inst_4.INIT_RAM_2F = 256'h4428290228502900150000280228155029001500000028022815442829286002;
defparam sp_inst_4.INIT_RAM_30 = 256'h0315002A150229024C0228032900150000280228155029001500000028022815;
defparam sp_inst_4.INIT_RAM_31 = 256'h4C022803290315150229024C02280329280028282829290229024C0228032900;
defparam sp_inst_4.INIT_RAM_32 = 256'h2A0315290028152815290229024C022800282950290240002828152929022902;
defparam sp_inst_4.INIT_RAM_33 = 256'h025347290228030303035029031429031528150229024C022803290003031500;
defparam sp_inst_4.INIT_RAM_34 = 256'h022828035703150257021C02021C022929024C02282803572903152815022929;
defparam sp_inst_4.INIT_RAM_35 = 256'h150257021C02021C022929024C022828035703150257021C02021C022929024C;
defparam sp_inst_4.INIT_RAM_36 = 256'h021C022929024C022828035703150257021C02021C022929024C022828035703;
defparam sp_inst_4.INIT_RAM_37 = 256'h4C022828035703150257021C02021C022929024C022828035703150257021C02;
defparam sp_inst_4.INIT_RAM_38 = 256'h03150257021C02021C022929024C022828035703150257021C02021C02292902;
defparam sp_inst_4.INIT_RAM_39 = 256'h02021C022929024C022828035703150257021C02021C022929024C0228280357;
defparam sp_inst_4.INIT_RAM_3A = 256'h024C022828035703150257021C02021C022929024C022828035703150257021C;
defparam sp_inst_4.INIT_RAM_3B = 256'h5703151457021C02021C022929024C022828035703150357021C02021C022929;
defparam sp_inst_4.INIT_RAM_3C = 256'h1C02021C022929024C022828035703151457021C02021C022929024C02282803;
defparam sp_inst_4.INIT_RAM_3D = 256'h29024C022828035703151457021C02021C022929024C02282803570315145702;
defparam sp_inst_4.INIT_RAM_3E = 256'h035703151457021C02021C022929024C022828035703151457021C02021C0229;
defparam sp_inst_4.INIT_RAM_3F = 256'h021C02021C022929024C022828035703151457021C02021C022929024C022828;

SP sp_inst_5 (
    .DO({sp_inst_5_dout_w[15:0],sp_inst_5_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[11],ad[10]}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_5.READ_MODE = 1'b0;
defparam sp_inst_5.WRITE_MODE = 2'b01;
defparam sp_inst_5.BIT_WIDTH = 16;
defparam sp_inst_5.BLK_SEL = 3'b010;
defparam sp_inst_5.RESET_MODE = "SYNC";
defparam sp_inst_5.INIT_RAM_00 = 256'h02B21C0002802980298002BF4C00028028802880034057F80380157F140057F3;
defparam sp_inst_5.INIT_RAM_01 = 256'h2980298002BF4C00028028802880034057F80380157F140057F202A61C000281;
defparam sp_inst_5.INIT_RAM_02 = 256'h4C00028028802880034057F70380157F140057F202A51C00028102B11C000280;
defparam sp_inst_5.INIT_RAM_03 = 256'h2880034057F70380157F140057F202A31C00028102B01C0002802980298002BF;
defparam sp_inst_5.INIT_RAM_04 = 256'h0380157F140157F202A21C00028202AF1C0002802980298002BF4C0002802880;
defparam sp_inst_5.INIT_RAM_05 = 256'h57F102A11C00028202AF1C0002802980298002BF4C00028028802880034057F7;
defparam sp_inst_5.INIT_RAM_06 = 256'h028202AE1C0002802980298002BF4C00028028802880034057F70380157F1402;
defparam sp_inst_5.INIT_RAM_07 = 256'h02802980298002BF4C00028028802880034057F60380157F140457F102A01C00;
defparam sp_inst_5.INIT_RAM_08 = 256'h02BF4C00028028802880034057F60380157F140857F1029F1C00028202AD1C00;
defparam sp_inst_5.INIT_RAM_09 = 256'h28802880034057F60380157F141057F0029D1C00028202AC1C00028029802980;
defparam sp_inst_5.INIT_RAM_0A = 256'h57F50380157F142057F0029C1C00028202AB1C0002802980298002BF4C000280;
defparam sp_inst_5.INIT_RAM_0B = 256'h144057F0029B1C00028202AB1C0002802980298002BF4C000280288028800340;
defparam sp_inst_5.INIT_RAM_0C = 256'h1C00028202AA1C0002802980298002BF4C00028028802880034057F50380157F;
defparam sp_inst_5.INIT_RAM_0D = 256'h1C0002802980298002BF4C00028028802880034057F50380157F148057EF029A;
defparam sp_inst_5.INIT_RAM_0E = 256'h298002BF4C00028028802880034057F40380157F150057EF02991C00028202A9;
defparam sp_inst_5.INIT_RAM_0F = 256'h29BF28800380157F57EF02971C00028302A81C00298014020380157F02802980;
defparam sp_inst_5.INIT_RAM_10 = 256'h40000340001728BF28BF500029BF034029BF001428BF28BF29BF28800380157F;
defparam sp_inst_5.INIT_RAM_11 = 256'h2880288003406FFF028028BF29BF028028BF4C0028800010004028BF02941C00;
defparam sp_inst_5.INIT_RAM_12 = 256'h034057F429BF28800380157F298014000380157F02802980298002BF4C000280;
defparam sp_inst_5.INIT_RAM_13 = 256'h157F297F037F006F004428800380157F02802980298002BF4C00028028802880;
defparam sp_inst_5.INIT_RAM_14 = 256'h1C0000152A7F298002800380157F298014000380157F293F0340006728800380;
defparam sp_inst_5.INIT_RAM_15 = 256'h0380157F298014000380157F0280298002BF4C00028028802880034057ED0293;
defparam sp_inst_5.INIT_RAM_16 = 256'h29BF0340004428800380157F02802980298002BF4C00028028800340293F2A00;
defparam sp_inst_5.INIT_RAM_17 = 256'h001002921C00004028BF6800028028BF2980001414010380157F28800380157F;
defparam sp_inst_5.INIT_RAM_18 = 256'h157F28800380157F57ED02911C00500029800380157F57ED02901C004C002880;
defparam sp_inst_5.INIT_RAM_19 = 256'h02802980298002BF4C000280288028800340034050002980001403BF15FF0380;
defparam sp_inst_5.INIT_RAM_1A = 256'h00670240288002A51CC74000001557F20284400003402A3F293F2A000380157F;
defparam sp_inst_5.INIT_RAM_1B = 256'h57F3400003402A3F57F2028457F002800015288002A41CC7298002A41CC70015;
defparam sp_inst_5.INIT_RAM_1C = 256'h028029800280157F5C00028028BF29BF2880157F5000293F28800380157F29BF;
defparam sp_inst_5.INIT_RAM_1D = 256'h293F28800380157F298028BF157F500029800280157F29BF400028BF500029BF;
defparam sp_inst_5.INIT_RAM_1E = 256'h28800340290002BF0380157F290002800380157F400003402A3F43FF0340283F;
defparam sp_inst_5.INIT_RAM_1F = 256'h028028802880034057EF57EB028A1C0057EF02802980298002BF4C0002802880;
defparam sp_inst_5.INIT_RAM_20 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C004C00;
defparam sp_inst_5.INIT_RAM_21 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_22 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_23 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_24 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_25 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_26 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_27 = 256'h2E2E2E2E2E2E00000A0D20203A636620203A696C3C201C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_28 = 256'h2E2E000078253A6C6E617965746E63752D2D00002E2E2E2E2E2E2E2E495F4F53;
defparam sp_inst_5.INIT_RAM_29 = 256'h2E2E2E2E2E2E44412E2E2E2E2E2E00002E2E2E2E2E2E2E2E414641422E2E2E2E;
defparam sp_inst_5.INIT_RAM_2A = 256'h1C001C001C001C001C001C0000002E2E7572746E726163206D69657200000A2E;
defparam sp_inst_5.INIT_RAM_2B = 256'h646E5F715F30697069741C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_2C = 256'h5F33697069740072646E5F715F32697069740072646E5F715F31697069740072;
defparam sp_inst_5.INIT_RAM_2D = 256'h69740072646E5F715F35697069740072646E5F715F34697069740072646E5F71;
defparam sp_inst_5.INIT_RAM_2E = 256'h646E5F715F30697069740072646E5F715F37697069740072646E5F715F366970;
defparam sp_inst_5.INIT_RAM_2F = 256'h5F33697069740072646E5F715F32697069740072646E5F715F31697069740072;
defparam sp_inst_5.INIT_RAM_30 = 256'h69740072646E5F715F35697069740072646E5F715F34697069740072646E5F71;
defparam sp_inst_5.INIT_RAM_31 = 256'h646E5F715F30697069740072646E5F715F37697069740072646E5F715F366970;
defparam sp_inst_5.INIT_RAM_32 = 256'h5F33697069740072646E5F715F32697069740072646E5F715F31697069740072;
defparam sp_inst_5.INIT_RAM_33 = 256'h69740072646E5F715F35697069740072646E5F715F34697069740072646E5F71;
defparam sp_inst_5.INIT_RAM_34 = 256'h646E5F715F30697069740072646E5F715F37697069740072646E5F715F366970;
defparam sp_inst_5.INIT_RAM_35 = 256'h5F33697069740072646E5F715F32697069740072646E5F715F31697069740072;
defparam sp_inst_5.INIT_RAM_36 = 256'h69740072646E5F715F35697069740072646E5F715F34697069740072646E5F71;
defparam sp_inst_5.INIT_RAM_37 = 256'h000000000072646E5F740072646E5F715F37697069740072646E5F715F366970;

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(sp_inst_0_dout[0]),
  .I1(sp_inst_2_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[1]),
  .I0(sp_inst_0_dout[1]),
  .I1(sp_inst_2_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(dout[2]),
  .I0(sp_inst_0_dout[2]),
  .I1(sp_inst_2_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(dout[3]),
  .I0(sp_inst_0_dout[3]),
  .I1(sp_inst_2_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[4]),
  .I0(sp_inst_0_dout[4]),
  .I1(sp_inst_2_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(dout[5]),
  .I0(sp_inst_0_dout[5]),
  .I1(sp_inst_2_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(dout[6]),
  .I0(sp_inst_0_dout[6]),
  .I1(sp_inst_2_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_23 (
  .O(dout[7]),
  .I0(sp_inst_0_dout[7]),
  .I1(sp_inst_2_dout[7]),
  .S0(dff_q_0)
);
MUX2 mux_inst_26 (
  .O(dout[8]),
  .I0(sp_inst_1_dout[8]),
  .I1(sp_inst_2_dout[8]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(dout[9]),
  .I0(sp_inst_1_dout[9]),
  .I1(sp_inst_2_dout[9]),
  .S0(dff_q_0)
);
MUX2 mux_inst_32 (
  .O(dout[10]),
  .I0(sp_inst_1_dout[10]),
  .I1(sp_inst_2_dout[10]),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(dout[11]),
  .I0(sp_inst_1_dout[11]),
  .I1(sp_inst_2_dout[11]),
  .S0(dff_q_0)
);
MUX2 mux_inst_38 (
  .O(dout[12]),
  .I0(sp_inst_1_dout[12]),
  .I1(sp_inst_2_dout[12]),
  .S0(dff_q_0)
);
MUX2 mux_inst_41 (
  .O(dout[13]),
  .I0(sp_inst_1_dout[13]),
  .I1(sp_inst_2_dout[13]),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(dout[14]),
  .I0(sp_inst_1_dout[14]),
  .I1(sp_inst_2_dout[14]),
  .S0(dff_q_0)
);
MUX2 mux_inst_47 (
  .O(dout[15]),
  .I0(sp_inst_1_dout[15]),
  .I1(sp_inst_2_dout[15]),
  .S0(dff_q_0)
);
MUX2 mux_inst_50 (
  .O(dout[16]),
  .I0(sp_inst_3_dout[16]),
  .I1(sp_inst_5_dout[16]),
  .S0(dff_q_0)
);
MUX2 mux_inst_53 (
  .O(dout[17]),
  .I0(sp_inst_3_dout[17]),
  .I1(sp_inst_5_dout[17]),
  .S0(dff_q_0)
);
MUX2 mux_inst_56 (
  .O(dout[18]),
  .I0(sp_inst_3_dout[18]),
  .I1(sp_inst_5_dout[18]),
  .S0(dff_q_0)
);
MUX2 mux_inst_59 (
  .O(dout[19]),
  .I0(sp_inst_3_dout[19]),
  .I1(sp_inst_5_dout[19]),
  .S0(dff_q_0)
);
MUX2 mux_inst_62 (
  .O(dout[20]),
  .I0(sp_inst_3_dout[20]),
  .I1(sp_inst_5_dout[20]),
  .S0(dff_q_0)
);
MUX2 mux_inst_65 (
  .O(dout[21]),
  .I0(sp_inst_3_dout[21]),
  .I1(sp_inst_5_dout[21]),
  .S0(dff_q_0)
);
MUX2 mux_inst_68 (
  .O(dout[22]),
  .I0(sp_inst_3_dout[22]),
  .I1(sp_inst_5_dout[22]),
  .S0(dff_q_0)
);
MUX2 mux_inst_71 (
  .O(dout[23]),
  .I0(sp_inst_3_dout[23]),
  .I1(sp_inst_5_dout[23]),
  .S0(dff_q_0)
);
MUX2 mux_inst_74 (
  .O(dout[24]),
  .I0(sp_inst_4_dout[24]),
  .I1(sp_inst_5_dout[24]),
  .S0(dff_q_0)
);
MUX2 mux_inst_77 (
  .O(dout[25]),
  .I0(sp_inst_4_dout[25]),
  .I1(sp_inst_5_dout[25]),
  .S0(dff_q_0)
);
MUX2 mux_inst_80 (
  .O(dout[26]),
  .I0(sp_inst_4_dout[26]),
  .I1(sp_inst_5_dout[26]),
  .S0(dff_q_0)
);
MUX2 mux_inst_83 (
  .O(dout[27]),
  .I0(sp_inst_4_dout[27]),
  .I1(sp_inst_5_dout[27]),
  .S0(dff_q_0)
);
MUX2 mux_inst_86 (
  .O(dout[28]),
  .I0(sp_inst_4_dout[28]),
  .I1(sp_inst_5_dout[28]),
  .S0(dff_q_0)
);
MUX2 mux_inst_89 (
  .O(dout[29]),
  .I0(sp_inst_4_dout[29]),
  .I1(sp_inst_5_dout[29]),
  .S0(dff_q_0)
);
MUX2 mux_inst_92 (
  .O(dout[30]),
  .I0(sp_inst_4_dout[30]),
  .I1(sp_inst_5_dout[30]),
  .S0(dff_q_0)
);
MUX2 mux_inst_95 (
  .O(dout[31]),
  .I0(sp_inst_4_dout[31]),
  .I1(sp_inst_5_dout[31]),
  .S0(dff_q_0)
);
endmodule //Gowin_SP_Instr
