//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Sat Mar 02 01:16:40 2024

module Gowin_SP_Instr (dout, clk, oce, ce, reset, wre, ad, din);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [11:0] ad;
input [31:0] din;

wire [23:0] sp_inst_0_dout_w;
wire [7:0] sp_inst_0_dout;
wire [23:0] sp_inst_1_dout_w;
wire [15:8] sp_inst_1_dout;
wire [15:0] sp_inst_2_dout_w;
wire [15:0] sp_inst_2_dout;
wire [23:0] sp_inst_3_dout_w;
wire [23:16] sp_inst_3_dout;
wire [23:0] sp_inst_4_dout_w;
wire [31:24] sp_inst_4_dout;
wire [15:0] sp_inst_5_dout_w;
wire [31:16] sp_inst_5_dout;
wire dff_q_0;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],sp_inst_0_dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b01;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h8CEC8C8C2C2C0C2C2CAC8C80ACAD0D8C0CCF8EEF2F8C2CAD0F900FF0EF4F000D;
defparam sp_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000200020006323800C2C8C6C2C;
defparam sp_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_20 = 256'hA08DA08DA08DA08DA08D0CA3A1ABAAA9A8A7A6A5A4B4B3B2B1B0AFAEADAC5535;
defparam sp_inst_0.INIT_RAM_21 = 256'hA5A4B4B3B2B1B0AFAEADAC550000A08D000000000000000000000000A08DA08D;
defparam sp_inst_0.INIT_RAM_22 = 256'hC6C5C4767661632063766100000485CCCC8C767661630015A3A1ABAAA9A8A7A6;
defparam sp_inst_0.INIT_RAM_23 = 256'hCCCC07A0CCCECDACCDCECDCC0780AECDCC00C0CCCC00FF04CC0CCC80CC80CCC7;
defparam sp_inst_0.INIT_RAM_24 = 256'h008C8C8CCC8D0CCDCC0C008CACCD8CCC8DCCCD00CCCC8CCEADCECDCC9FCCCC8C;
defparam sp_inst_0.INIT_RAM_25 = 256'hCCFF84CCFF04AC0CCD00C47676616320637661840C0CCCCC8CCCFF848C8C8CCC;
defparam sp_inst_0.INIT_RAM_26 = 256'h00C0CCCCCC8CCCCBCAC9C8C7C6C5C47676616320637661840C9FCCCC8CCCCC8C;
defparam sp_inst_0.INIT_RAM_27 = 256'hCCCC8CCCFF848CCC808CAC8C2C8DAC0D8C8CACCD8CCCCC0CAC0CCDCC8CACCDCC;
defparam sp_inst_0.INIT_RAM_28 = 256'h078CCC00CC8CCCCC8CCCFF84C506078CCC00CC8CCCCC8CCCFF848C8CCC00CC8C;
defparam sp_inst_0.INIT_RAM_29 = 256'hFF84C506078CCC00CC8CCCCC8CCCFF84C506078CCC00CC8CCCCC8CCCFF84C506;
defparam sp_inst_0.INIT_RAM_2A = 256'h00C0CC8CCC00CC8CCCFF0400CC8CCCCC8CCCFF84C506078CCC00CC8CCCCC8CCC;
defparam sp_inst_0.INIT_RAM_2B = 256'hCD00C0FF8D0C8DACCD8CCC8D0C8DACCD8CCCCC8CCCCCAC8C8CCCCE8CCCAD0CCD;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000FF04FF8D0C8DACCD8CCC8D0C8DACCD8CCCCC8CCCCCAC8C8CCCCE8CCCAD0C;
defparam sp_inst_0.INIT_RAM_2D = 256'h8C8CCC00CCACC476766320637661840C9F8CACCDCCCC8CCCFF84CCFF04AC0CCD;
defparam sp_inst_0.INIT_RAM_2E = 256'h002C0C7676632063760020767663206376008C0C767663206376008DCDCC9F8C;
defparam sp_inst_0.INIT_RAM_2F = 256'h767663206376008DADAD0C767663206376008DCCADCC8DCCC5C4767663206376;
defparam sp_inst_0.INIT_RAM_30 = 256'h8C0C8D8C8C0C8DCDCD0C8E0CC476766320637684CCC000CC0C80ACCC8D0CC0C4;
defparam sp_inst_0.INIT_RAM_31 = 256'hACC476766320637661000084C485CC8D0D8CCCCC8C76766163206376008DADAD;
defparam sp_inst_0.INIT_RAM_32 = 256'h8DCC8D8CCC8DCC8DCC8D8CCC80CCAC8CCC8DCC8DCC8D8CCC8DCD8CADCD8CCCCC;
defparam sp_inst_0.INIT_RAM_33 = 256'h766163008D0DCCCC2CFF767661632063760080CCAC8CCC8DCC8DCC8D8CCC8DCC;
defparam sp_inst_0.INIT_RAM_34 = 256'h6100FF840C05FF842405C626767661632063766100FF840C05FF842405C62676;
defparam sp_inst_0.INIT_RAM_35 = 256'hFF842405C626767661632063766100FF840C05FF842405C62676766163206376;
defparam sp_inst_0.INIT_RAM_36 = 256'h767661632063766100FF840C05FF842405C626767661632063766100FF840C05;
defparam sp_inst_0.INIT_RAM_37 = 256'h766100FF840C05FF842405C626767661632063766100FF840C05FF842405C626;
defparam sp_inst_0.INIT_RAM_38 = 256'h05FF842405C626767661632063766100FF840C05FF842405C626767661632063;
defparam sp_inst_0.INIT_RAM_39 = 256'h26767661632063766100FF840C05FF842405C626767661632063766100FF840C;
defparam sp_inst_0.INIT_RAM_3A = 256'h63766100FF840C05FF842405C626767661632063766100FF840C05FF842405C6;
defparam sp_inst_0.INIT_RAM_3B = 256'h0C45FF842405C626767661632063766100FF840C25FF842405C6267676616320;
defparam sp_inst_0.INIT_RAM_3C = 256'hC626767661632063766100FF840C85FF842405C626767661632063766100FF84;
defparam sp_inst_0.INIT_RAM_3D = 256'h2063766100FF840C05FF842405C626767661632063766100FF840C05FF842405;
defparam sp_inst_0.INIT_RAM_3E = 256'h840C05FF842405C626767661632063766100FF840C05FF842405C62676766163;
defparam sp_inst_0.INIT_RAM_3F = 256'h05C626767661632063766100FF840C05FF842405C626767661632063766100FF;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[23:0],sp_inst_1_dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:8]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b01;
defparam sp_inst_1.BIT_WIDTH = 8;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'hFDE311FD0010003000F911011101000100D135010001001102350235E1002000;
defparam sp_inst_1.INIT_RAM_01 = 256'h000000000000000000000000000000000000000000800028F00001204041A044;
defparam sp_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_20 = 256'h2D812D412D212D1165F114425262728292A2B2C2D2728292A2B2C2D2E2F200C4;
defparam sp_inst_1.INIT_RAM_21 = 256'hC2D2728292A2B2C2D2E2F20004640D0114581CC424AC2C7834F43CB42D012D01;
defparam sp_inst_1.INIT_RAM_22 = 256'h526272C0A0B04000806070008CD001BEBE008060708038C4425262728292A2B2;
defparam sp_inst_1.INIT_RAM_23 = 256'hB2920009359252C135C2B25D0009B1925250B292720C87B49230721D72254242;
defparam sp_inst_1.INIT_RAM_24 = 256'h1481C18182192482820008C131C2FDA21DB2A274A23135B531B2B262B192B205;
defparam sp_inst_1.INIT_RAM_25 = 256'h723301BE3F340D28BE3072C0A0B04000C0A0B001008CA2A2FDA29701815D8182;
defparam sp_inst_1.INIT_RAM_26 = 256'h30B2A272729182726252423222123200E0F08000C0A0B00100C5BEBE01727205;
defparam sp_inst_1.INIT_RAM_27 = 256'hB2A211A2DB0101A2010131F10089AD4C6D01313205B29204E5948E8E013132B2;
defparam sp_inst_1.INIT_RAM_28 = 256'h0401A230B205B2A211A2130192280001A268B205B2A211A20F018101A298B205;
defparam sp_inst_1.INIT_RAM_29 = 256'h6B0192080001A2C0B205B2A211A2A30192200001A2F8B205B2A211A2DB019228;
defparam sp_inst_1.INIT_RAM_2A = 256'h3C92B205B238B205B2D39450B205B2A211A2330192400001A288B205B2A211A2;
defparam sp_inst_1.INIT_RAM_2B = 256'h923C92BB95E401313205B2D9C001313205B2B205B292314101313205B2312892;
defparam sp_inst_1.INIT_RAM_2C = 256'h2400B7943F95E401313205B25DC001313205B2B205B292314101313205B23128;
defparam sp_inst_1.INIT_RAM_2D = 256'h8115B200AE00B28070800080E0F00100C5013132B2B205B28F018E9B340D288E;
defparam sp_inst_1.INIT_RAM_2E = 256'h0010044030C000403000044030C00040300001104030C00080700001AEB2F181;
defparam sp_inst_1.INIT_RAM_2F = 256'hC0B04000403000D1A9B4D64030C00080700031B231A231B2A2B2807080004030;
defparam sp_inst_1.INIT_RAM_30 = 256'h0DD481010DD40135B2DA01DAB280708000C0B001B2B208B20411B17201DAB272;
defparam sp_inst_1.INIT_RAM_31 = 256'h00B2807080008060700018E0FF01BE010431FFBE008060708000807000018105;
defparam sp_inst_1.INIT_RAM_32 = 256'h11B24511B241B241B20541B231B20D11B231B231B20531B201AE3531B201B2AE;
defparam sp_inst_1.INIT_RAM_33 = 256'h2030C0000104B2B2004F806070800080700021B20D11B221B221B20521B241B2;
defparam sp_inst_1.INIT_RAM_34 = 256'h30001B81D608D3F00060D000402030C000402030006781D6041F20004CA00040;
defparam sp_inst_1.INIT_RAM_35 = 256'h3B9000883000402030C00040203000CF81D61087C000740000402030C0004020;
defparam sp_inst_1.INIT_RAM_36 = 256'h402030C000402030003781D640EF60009C6000402030C000402030008381D620;
defparam sp_inst_1.INIT_RAM_37 = 256'h2030009F81D600570000C4C000402030C00040203000EB81D680A33000B09000;
defparam sp_inst_1.INIT_RAM_38 = 256'h00BFA000F02000402030C000402030005381D6000BD000DCF000402030C00040;
defparam sp_inst_1.INIT_RAM_39 = 256'h00402030C00040203000BB81D600737000085000402030C000402030000781D6;
defparam sp_inst_1.INIT_RAM_3A = 256'h402030002381D600DB100038B000402030C000402030006F81D6002740002080;
defparam sp_inst_1.INIT_RAM_3B = 256'hD60043B000601000402030C00040203000D781D6008FE0004CE000402030C000;
defparam sp_inst_1.INIT_RAM_3C = 256'h7000402030C000402030003F81D600F78000784000402030C000402030008B81;
defparam sp_inst_1.INIT_RAM_3D = 256'h0040203000A781D6025F2000ACA000402030C00040203000F381D601AB500090;
defparam sp_inst_1.INIT_RAM_3E = 256'h81D608C7C000DC0000402030C000402030005B81D60413F000C4D000402030C0;
defparam sp_inst_1.INIT_RAM_3F = 256'h0C6000402030C00040203000C381D6107B9000F43000402030C000402030000F;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[15:0],sp_inst_2_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[11],ad[10]}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b01;
defparam sp_inst_2.BIT_WIDTH = 16;
defparam sp_inst_2.BLK_SEL = 3'b010;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'h407620763061C0630020406320763061000077FF8184D60C20052FFF60840024;
defparam sp_inst_2.INIT_RAM_01 = 256'hC063002040632076306100002BFF8184D60C4005E3FF30840024200590C60026;
defparam sp_inst_2.INIT_RAM_02 = 256'h207630610000DFFF8184D60C800597FF008400243405C0C60026407620763061;
defparam sp_inst_2.INIT_RAM_03 = 256'h93FF8184D60C00054BFFD08400044C05F0C60026407620763061C06300204063;
defparam sp_inst_2.INIT_RAM_04 = 256'h0005FFFFA0840004640520C60026407620763061C06300204063207630610000;
defparam sp_inst_2.INIT_RAM_05 = 256'h00047C0550C60026407620763061C0630020406320763061000047FF8184D60C;
defparam sp_inst_2.INIT_RAM_06 = 256'h0026407620763061C06300204063207630610000FBFF8184D60C0005B3FF7084;
defparam sp_inst_2.INIT_RAM_07 = 256'h3061C06300204063207630610000AFFF8184D60C000567FF40840004940580C6;
defparam sp_inst_2.INIT_RAM_08 = 256'h406320763061000063FF8184D60C00051BFF10840004AC05B0C6002640762076;
defparam sp_inst_2.INIT_RAM_09 = 256'h000017FF8184D60C0005CFFFE0840004C405E0C60026407620763061C0630020;
defparam sp_inst_2.INIT_RAM_0A = 256'hD60C000583FFB0840004E00510C60026407620763061C0630020406320763061;
defparam sp_inst_2.INIT_RAM_0B = 256'h80840004F80540C60026407620763061C06300204063207630610000CBFF8184;
defparam sp_inst_2.INIT_RAM_0C = 256'h70C60026407620763061C063002040632076306100007FFF8184D60C000537FF;
defparam sp_inst_2.INIT_RAM_0D = 256'h6076706180630020406320763061000033FF8184D60C0005EBFF508400041005;
defparam sp_inst_2.INIT_RAM_0E = 256'hD60CA2CC318C818CD60C8FFFE0840004C00560C60026018D000DF18CD60C8076;
defparam sp_inst_2.INIT_RAM_0F = 256'h000D2180058CB1ACB2CCA2CD4000B2C00000A2CCB1AC92CCA2CD92CC018C818C;
defparam sp_inst_2.INIT_RAM_10 = 256'h8063607670610000BD8D7C0CB2CDB2CC058CB2CC0181018C31AC898CB2CCB1AD;
defparam sp_inst_2.INIT_RAM_11 = 256'h7061000057FFB2CC018C118CD60C018D020DF18CD60C80766076706180630020;
defparam sp_inst_2.INIT_RAM_12 = 256'h118CD68CBACCFD8C818CC18C018C118CD68C8076607670618063002080636076;
defparam sp_inst_2.INIT_RAM_13 = 256'hA08400040185BACC018D3C0D118CD68C018D040DF18CD60CB6CC3D8C818C018C;
defparam sp_inst_2.INIT_RAM_14 = 256'h018C098CD18C018D080DF18CD60C8076707680630020806360767061000037FF;
defparam sp_inst_2.INIT_RAM_15 = 256'hD60CB2CC7D8CCD8C018C118CD60C80766076706180630020806370760000BECC;
defparam sp_inst_2.INIT_RAM_16 = 256'h018C31ACE18C000C898DB2CC718D400CB2CD018DB5CDF00DF18CD60C018E118C;
defparam sp_inst_2.INIT_RAM_17 = 256'h118CD60C018E118CD60C4FFF208400043C000180118CD60C6BFFF08400040180;
defparam sp_inst_2.INIT_RAM_18 = 256'hD40C80766076706180630020806360767061000000000800018DB5CDFDADFEED;
defparam sp_inst_2.INIT_RAM_19 = 256'hBECCBFFF70840004D7FF00041980008C9BFF00042980058CBECCBECC018C158C;
defparam sp_inst_2.INIT_RAM_1A = 256'h218CBECC018D100D0D8CD40C93FF608400040185BACCBACC018CD10C3580118C;
defparam sp_inst_2.INIT_RAM_1B = 256'h0000018DFC0D0D8CD40C018D200D0D8CD40CC7FF0184B6CCB6CC018CD00C2D80;
defparam sp_inst_2.INIT_RAM_1C = 256'h2076306100001BFF0BFF908400044BFF407620763061C0630020806360767061;
defparam sp_inst_2.INIT_RAM_1D = 256'h15F415F4156C1670167016701670167016701670167016701670155400204063;
defparam sp_inst_2.INIT_RAM_1E = 256'h16701670167016701670167016701670167015F415F415F415F415F415F415F4;
defparam sp_inst_2.INIT_RAM_1F = 256'h1670167016701670167016701670167016701670167016701670167016701670;
defparam sp_inst_2.INIT_RAM_20 = 256'h14E4167016701670167016701670167016701670167016701670167016701670;
defparam sp_inst_2.INIT_RAM_21 = 256'h16701670151C14AC16701670167016701670167016701670167016701474140C;
defparam sp_inst_2.INIT_RAM_22 = 256'h2E2E2E0A00003E2073256E756425656E20200A0D151C16701670143C167013E0;
defparam sp_inst_2.INIT_RAM_23 = 256'h000A7830656E68434B3A49686F742D0A0D0A2E2E2E2E2E2E544E54462E2E2E2E;
defparam sp_inst_2.INIT_RAM_24 = 256'h2E2E2E432E2E2E2E2E2E2E0A0D0A2E2E2E2E2E2E4C495F542E2E2E2E2E2E2E0A;
defparam sp_inst_2.INIT_RAM_25 = 256'h76632031617500002E7472726E696165207269546C6168706550000D2E2E2E2E;
defparam sp_inst_2.INIT_RAM_26 = 256'h1B701B241AD81A8C1A4019F4000A747072656920656C726554206F4300002578;
defparam sp_inst_2.INIT_RAM_27 = 256'h20301FE41F981F4C1F001EB41E681E1C1DD01D841D381CEC1CA01C541C081BBC;
defparam sp_inst_2.INIT_RAM_28 = 256'h261426142614261425C42614232822DC2290224421F821AC2160211420C8207C;
defparam sp_inst_2.INIT_RAM_29 = 256'h61687269616F675F786525E02614261426142614261426142614261426142614;
defparam sp_inst_2.INIT_RAM_2A = 256'h616F675F7865656C61687269616F675F7865656C61687269616F675F7865656C;
defparam sp_inst_2.INIT_RAM_2B = 256'h7865656C61687269616F675F7865656C61687269616F675F7865656C61687269;
defparam sp_inst_2.INIT_RAM_2C = 256'h61687269626F675F7865656C61687269616F675F7865656C61687269616F675F;
defparam sp_inst_2.INIT_RAM_2D = 256'h626F675F7865656C61687269626F675F7865656C61687269626F675F7865656C;
defparam sp_inst_2.INIT_RAM_2E = 256'h7865656C61687269626F675F7865656C61687269626F675F7865656C61687269;
defparam sp_inst_2.INIT_RAM_2F = 256'h61687269636F675F7865656C61687269626F675F7865656C61687269626F675F;
defparam sp_inst_2.INIT_RAM_30 = 256'h636F675F7865656C61687269636F675F7865656C61687269636F675F7865656C;
defparam sp_inst_2.INIT_RAM_31 = 256'h7865656C61687269636F675F7865656C61687269636F675F7865656C61687269;
defparam sp_inst_2.INIT_RAM_32 = 256'h61687269646F675F7865656C61687269636F675F7865656C61687269636F675F;
defparam sp_inst_2.INIT_RAM_33 = 256'h646F675F7865656C61687269646F675F7865656C61687269646F675F7865656C;
defparam sp_inst_2.INIT_RAM_34 = 256'h7865656C61687269646F675F7865656C61687269646F675F7865656C61687269;
defparam sp_inst_2.INIT_RAM_35 = 256'h00000000656C61687865656C61687269646F675F7865656C61687269646F675F;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[23:0],sp_inst_3_dout[23:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[23:16]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b01;
defparam sp_inst_3.BIT_WIDTH = 8;
defparam sp_inst_3.BLK_SEL = 3'b000;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'hBFFF00BF0000150038FF80800080008000FF10800080008080108010B5380015;
defparam sp_inst_3.INIT_RAM_01 = 256'h000000000000000000000000000000000000000000480019BD0000800688EC06;
defparam sp_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_20 = 256'h0040004000400040006E00BEBEBEBEBEBEBEBEBEBEBFBFBFBFBFBFBFBFBF0000;
defparam sp_inst_3.INIT_RAM_21 = 256'hBEBEBFBFBFBFBFBFBFBFBF000015004100160012001400140013001300600042;
defparam sp_inst_3.INIT_RAM_22 = 256'hBEBEBE818181BE0080808040057F153F3F15808080BF4800BEBEBEBEBEBEBEBE;
defparam sp_inst_3.INIT_RAM_23 = 256'hBFBF2A0021BFBE3E10BFBF002A0021BFBE00BFBFBE00FF80BF11BE00BE00BEBE;
defparam sp_inst_3.INIT_RAM_24 = 256'h00678067BF0080BFBF15003E10BFBFBF00BFBF00BF15131312BFBFBEFFBFBF80;
defparam sp_inst_3.INIT_RAM_25 = 256'hBFFE153FFE8000803F00BF808080BF008181811515FFBFBFBFBFFE15678167BF;
defparam sp_inst_3.INIT_RAM_26 = 256'h03BFBFBFBFBF8080808080808080BF818080BE008080801515FF3F3F00BFBF80;
defparam sp_inst_3.INIT_RAM_27 = 256'hBFBF80BFFE1580BF0080108D00400281BF0010BF80BFBF8002803F3F0010BFBF;
defparam sp_inst_3.INIT_RAM_28 = 256'h8080BF02BF80BFBF80BFFD15BF801580BF02BF80BFBF80BFFD156780BF02BF80;
defparam sp_inst_3.INIT_RAM_29 = 256'hFC15BF801580BF01BF80BFBF80BFFC15BF801580BF01BF80BFBF80BFFC15BF80;
defparam sp_inst_3.INIT_RAM_2A = 256'h00BFBF80BF01BF80BFFB8001BF80BFBF80BFFC15BF801580BF01BF80BFBF80BF;
defparam sp_inst_3.INIT_RAM_2B = 256'hBF00BFFDFF800010BF80BFFD800010BF80BFBF80BFBF10BF0010BF80BF1C80BF;
defparam sp_inst_3.INIT_RAM_2C = 256'h0040FA80FDFF800010BF80BFFD800010BF80BFBF80BFBF10BF0010BF80BF1C80;
defparam sp_inst_3.INIT_RAM_2D = 256'h6700BF403F15BF8080BF008180801515FC0010BFBFBF80BFFA153FFA8000803F;
defparam sp_inst_3.INIT_RAM_2E = 256'h4001808080BF00808040018080BF0080804000808080BF00808040003FBFFF40;
defparam sp_inst_3.INIT_RAM_2F = 256'h8080BF0080804080964A7F8080BF0080804080BF15BF80BFBFBF8080BF008080;
defparam sp_inst_3.INIT_RAM_30 = 256'h807F6700807F8015BF7F807FBF8080BF00808015BFBF00BF800014BF807FBFBF;
defparam sp_inst_3.INIT_RAM_31 = 256'h15BF8080BF0080808040009CC7153F80809DC73F15808080BF00808040006780;
defparam sp_inst_3.INIT_RAM_32 = 256'h80BF0080BF80BF80BF8080BF80BF0080BF80BF80BF8080BF003F1080BF80BF3F;
defparam sp_inst_3.INIT_RAM_33 = 256'h8080BF008080BFBF00FD808080BF0080804080BF0080BF80BF80BF8080BF80BF;
defparam sp_inst_3.INIT_RAM_34 = 256'h8040FD807F80F8B800808000808080BF0080808040FD807F80F9BA0080810080;
defparam sp_inst_3.INIT_RAM_35 = 256'hF8B60080BF00808080BF0080808040FC807F80F8B700808000808080BF008080;
defparam sp_inst_3.INIT_RAM_36 = 256'h808080BF0080808040FC807F80F7B50080BE00808080BF0080808040FC807F80;
defparam sp_inst_3.INIT_RAM_37 = 256'h808040FB807F81F7B30080BC00808080BF0080808040FB807F80F7B40080BD00;
defparam sp_inst_3.INIT_RAM_38 = 256'h84F6B00080BB00808080BF0080808040FB807F82F7B10080BB00808080BF0080;
defparam sp_inst_3.INIT_RAM_39 = 256'h00808080BF0080808040FA807F88F6AF0081BA00808080BF0080808040FB807F;
defparam sp_inst_3.INIT_RAM_3A = 256'h80808040FA807FA0F5AD0081B800808080BF0080808040FA807F90F6AE0081B9;
defparam sp_inst_3.INIT_RAM_3B = 256'h7F00F5AA0081B700808080BF0080808040F9807F00F5AB0081B700808080BF00;
defparam sp_inst_3.INIT_RAM_3C = 256'hB500808080BF0080808040F9807F00F4A90081B600808080BF0080808040F980;
defparam sp_inst_3.INIT_RAM_3D = 256'h0080808040F8807F00F4A70081B400808080BF0080808040F8807F00F4A80081;
defparam sp_inst_3.INIT_RAM_3E = 256'h807F00F3A40081B300808080BF0080808040F8807F00F4A50081B300808080BF;
defparam sp_inst_3.INIT_RAM_3F = 256'h82B100808080BF0080808040F7807F00F3A30081B200808080BF0080808040F8;

SP sp_inst_4 (
    .DO({sp_inst_4_dout_w[23:0],sp_inst_4_dout[31:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:24]})
);

defparam sp_inst_4.READ_MODE = 1'b0;
defparam sp_inst_4.WRITE_MODE = 2'b01;
defparam sp_inst_4.BIT_WIDTH = 8;
defparam sp_inst_4.BLK_SEL = 3'b000;
defparam sp_inst_4.RESET_MODE = "SYNC";
defparam sp_inst_4.INIT_RAM_00 = 256'h0315040314040004145F022958031503155F0003150315022900280003145000;
defparam sp_inst_4.INIT_RAM_01 = 256'h00000000000000000000000000000000000000004C064C540315040304031404;
defparam sp_inst_4.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_20 = 256'h4403440344034403400304292929292929292929292929292929292929291504;
defparam sp_inst_4.INIT_RAM_21 = 256'h2828282828282828282828155054400350545054505450545054505444034403;
defparam sp_inst_4.INIT_RAM_22 = 256'h292929022929024C022828035415002A29000229290206042828282828282828;
defparam sp_inst_4.INIT_RAM_23 = 256'h2829005C0028282900022800005C002828502929285057022900286428402829;
defparam sp_inst_4.INIT_RAM_24 = 256'h5000020028600228290050280002022860282850290000000028282847282902;
defparam sp_inst_4.INIT_RAM_25 = 256'h2857002A57025C02285029022929024C02282800006328290228570000020028;
defparam sp_inst_4.INIT_RAM_26 = 256'h502929282902022929292929292929022929024C02282800004728292A282902;
defparam sp_inst_4.INIT_RAM_27 = 256'h28290228570028284C2800021C00680202280028022829025C0228292A002828;
defparam sp_inst_4.INIT_RAM_28 = 256'h0228285029022829022857002802002828502902282902285700002828502902;
defparam sp_inst_4.INIT_RAM_29 = 256'h5700280200282850290228290228570028020028285029022829022857002802;
defparam sp_inst_4.INIT_RAM_2A = 256'h5029290228502902285702502902282902285700280200282850290228290228;
defparam sp_inst_4.INIT_RAM_2B = 256'h2850295367022800280228670228002802282902282900022800280228000228;
defparam sp_inst_4.INIT_RAM_2C = 256'h5003570253670228002802286702280028022829022829000228002802280002;
defparam sp_inst_4.INIT_RAM_2D = 256'h002A28032900290229024C0228280000472800282829022857002A57025C0228;
defparam sp_inst_4.INIT_RAM_2E = 256'h0304030229024C022803040229024C02280304030229024C022803292A284303;
defparam sp_inst_4.INIT_RAM_2F = 256'h0229024C022803290315150229024C02280329280028282829290229024C0228;
defparam sp_inst_4.INIT_RAM_30 = 256'h0315002A0315290028152815290229024C022800282950290240002828152929;
defparam sp_inst_4.INIT_RAM_31 = 256'h00290229024C0228280354021C002A2902021C2900022929024C022803290003;
defparam sp_inst_4.INIT_RAM_32 = 256'h282864282828282928022828292860282828282928022828292A002828282829;
defparam sp_inst_4.INIT_RAM_33 = 256'h29290250290228291557022929024C0228032928602828282829280228282928;
defparam sp_inst_4.INIT_RAM_34 = 256'h28035703150257021C02021C022929024C022828035703150257021C02021C02;
defparam sp_inst_4.INIT_RAM_35 = 256'h57021C02021C022929024C022828035703150257021C02021C022929024C0228;
defparam sp_inst_4.INIT_RAM_36 = 256'h022929024C022828035703150257021C02021C022929024C0228280357031502;
defparam sp_inst_4.INIT_RAM_37 = 256'h2828035703150257021C02021C022929024C022828035703150257021C02021C;
defparam sp_inst_4.INIT_RAM_38 = 256'h0257021C02021C022929024C022828035703150257021C02021C022929024C02;
defparam sp_inst_4.INIT_RAM_39 = 256'h1C022929024C022828035703150257021C02021C022929024C02282803570315;
defparam sp_inst_4.INIT_RAM_3A = 256'h022828035703150357021C02021C022929024C022828035703150257021C0202;
defparam sp_inst_4.INIT_RAM_3B = 256'h151457021C02021C022929024C022828035703151457021C02021C022929024C;
defparam sp_inst_4.INIT_RAM_3C = 256'h021C022929024C022828035703151457021C02021C022929024C022828035703;
defparam sp_inst_4.INIT_RAM_3D = 256'h4C022828035703151457021C02021C022929024C022828035703151457021C02;
defparam sp_inst_4.INIT_RAM_3E = 256'h03151457021C02021C022929024C022828035703151457021C02021C02292902;
defparam sp_inst_4.INIT_RAM_3F = 256'h02021C022929024C022828035703151457021C02021C022929024C0228280357;

SP sp_inst_5 (
    .DO({sp_inst_5_dout_w[15:0],sp_inst_5_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[11],ad[10]}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_5.READ_MODE = 1'b0;
defparam sp_inst_5.WRITE_MODE = 2'b01;
defparam sp_inst_5.BIT_WIDTH = 16;
defparam sp_inst_5.BLK_SEL = 3'b010;
defparam sp_inst_5.RESET_MODE = "SYNC";
defparam sp_inst_5.INIT_RAM_00 = 256'h02802980298002BF4C00028028802880034057F70380157F140057F302A21C00;
defparam sp_inst_5.INIT_RAM_01 = 256'h02BF4C00028028802880034057F70380157F140057F202A11C00028202B01C00;
defparam sp_inst_5.INIT_RAM_02 = 256'h28802880034057F60380157F140057F202A01C00028202AF1C00028029802980;
defparam sp_inst_5.INIT_RAM_03 = 256'h57F60380157F140157F2029E1C00028202AE1C0002802980298002BF4C000280;
defparam sp_inst_5.INIT_RAM_04 = 256'h140257F1029D1C00028202AE1C0002802980298002BF4C000280288028800340;
defparam sp_inst_5.INIT_RAM_05 = 256'h1C00028202AD1C0002802980298002BF4C00028028802880034057F60380157F;
defparam sp_inst_5.INIT_RAM_06 = 256'h1C0002802980298002BF4C00028028802880034057F50380157F140457F1029C;
defparam sp_inst_5.INIT_RAM_07 = 256'h298002BF4C00028028802880034057F50380157F140857F1029B1C00028202AC;
defparam sp_inst_5.INIT_RAM_08 = 256'h028028802880034057F50380157F141057F1029A1C00028202AB1C0002802980;
defparam sp_inst_5.INIT_RAM_09 = 256'h034057F50380157F142057F002981C00028202AA1C0002802980298002BF4C00;
defparam sp_inst_5.INIT_RAM_0A = 256'h157F144057F002971C00028202AA1C0002802980298002BF4C00028028802880;
defparam sp_inst_5.INIT_RAM_0B = 256'h02961C00028202A91C0002802980298002BF4C00028028802880034057F40380;
defparam sp_inst_5.INIT_RAM_0C = 256'h02A81C0002802980298002BF4C00028028802880034057F40380157F148057F0;
defparam sp_inst_5.INIT_RAM_0D = 256'h2980298002BF4C00028028802880034057F40380157F150057EF02951C000283;
defparam sp_inst_5.INIT_RAM_0E = 256'h157F29BF28800380157F57EF02931C00028302A71C00298014020380157F0280;
defparam sp_inst_5.INIT_RAM_0F = 256'h1C0040000340001728BF28BF500029BF034029BF001428BF28BF29BF28800380;
defparam sp_inst_5.INIT_RAM_10 = 256'h02802880288003406FFF028028BF29BF028028BF4C0028800010004028BF0296;
defparam sp_inst_5.INIT_RAM_11 = 256'h2880034057F329BF28800380157F298014000380157F02802980298002BF4C00;
defparam sp_inst_5.INIT_RAM_12 = 256'h0380157F297F037F006F004428800380157F02802980298002BF4C0002802880;
defparam sp_inst_5.INIT_RAM_13 = 256'h028F1C0000152A7F298002800380157F298014000380157F293F034000672880;
defparam sp_inst_5.INIT_RAM_14 = 256'h2A000380157F298014000380157F0280298002BF4C00028028802880034057EE;
defparam sp_inst_5.INIT_RAM_15 = 256'h157F29BF0340004428800380157F02802980298002BF4C00028028800340293F;
defparam sp_inst_5.INIT_RAM_16 = 256'h2880001002911C00004028BF6800028028BF2980001414010380157F28800380;
defparam sp_inst_5.INIT_RAM_17 = 256'h0380157F28800380157F57ED028D1C00500029800380157F57ED028C1C004C00;
defparam sp_inst_5.INIT_RAM_18 = 256'h157F02802980298002BF4C000280288028800340034050002980001403BF15FF;
defparam sp_inst_5.INIT_RAM_19 = 256'h2A3F57EC028B1C0057F102844000001557F10284400003402A3F293F2A000380;
defparam sp_inst_5.INIT_RAM_1A = 256'h03402A3F290002800380157F57EC028B1C0000152A3F293F2A00157F40000340;
defparam sp_inst_5.INIT_RAM_1B = 256'h0340290002BF0380157F290002800380157F57F100152A3F293F2A00157F4000;
defparam sp_inst_5.INIT_RAM_1C = 256'h28802880034057F057EC02891C0057F002802980298002BF4C00028028802880;
defparam sp_inst_5.INIT_RAM_1D = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C004C000280;
defparam sp_inst_5.INIT_RAM_1E = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_1F = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_20 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_21 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_22 = 256'h2E2E2E2E00000A0D20203A636620203A696C3C201C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_23 = 256'h000078253A6C6E617965746E63752D2D00002E2E2E2E2E2E2E2E495F4F532E2E;
defparam sp_inst_5.INIT_RAM_24 = 256'h2E2E2E2E44412E2E2E2E2E2E00002E2E2E2E2E2E2E2E414641422E2E2E2E2E2E;
defparam sp_inst_5.INIT_RAM_25 = 256'h303A6572747200000A2E7075657420726C63656D20737265697200000A2E2E2E;
defparam sp_inst_5.INIT_RAM_26 = 256'h1C001C001C001C001C001C0000002E2E7572746E726163206D69657200000A78;
defparam sp_inst_5.INIT_RAM_27 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_28 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_29 = 256'h646E5F715F30697069741C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_5.INIT_RAM_2A = 256'h5F33697069740072646E5F715F32697069740072646E5F715F31697069740072;
defparam sp_inst_5.INIT_RAM_2B = 256'h69740072646E5F715F35697069740072646E5F715F34697069740072646E5F71;
defparam sp_inst_5.INIT_RAM_2C = 256'h646E5F715F30697069740072646E5F715F37697069740072646E5F715F366970;
defparam sp_inst_5.INIT_RAM_2D = 256'h5F33697069740072646E5F715F32697069740072646E5F715F31697069740072;
defparam sp_inst_5.INIT_RAM_2E = 256'h69740072646E5F715F35697069740072646E5F715F34697069740072646E5F71;
defparam sp_inst_5.INIT_RAM_2F = 256'h646E5F715F30697069740072646E5F715F37697069740072646E5F715F366970;
defparam sp_inst_5.INIT_RAM_30 = 256'h5F33697069740072646E5F715F32697069740072646E5F715F31697069740072;
defparam sp_inst_5.INIT_RAM_31 = 256'h69740072646E5F715F35697069740072646E5F715F34697069740072646E5F71;
defparam sp_inst_5.INIT_RAM_32 = 256'h646E5F715F30697069740072646E5F715F37697069740072646E5F715F366970;
defparam sp_inst_5.INIT_RAM_33 = 256'h5F33697069740072646E5F715F32697069740072646E5F715F31697069740072;
defparam sp_inst_5.INIT_RAM_34 = 256'h69740072646E5F715F35697069740072646E5F715F34697069740072646E5F71;
defparam sp_inst_5.INIT_RAM_35 = 256'h000000000072646E5F740072646E5F715F37697069740072646E5F715F366970;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(sp_inst_0_dout[0]),
  .I1(sp_inst_2_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[1]),
  .I0(sp_inst_0_dout[1]),
  .I1(sp_inst_2_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(dout[2]),
  .I0(sp_inst_0_dout[2]),
  .I1(sp_inst_2_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(dout[3]),
  .I0(sp_inst_0_dout[3]),
  .I1(sp_inst_2_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[4]),
  .I0(sp_inst_0_dout[4]),
  .I1(sp_inst_2_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(dout[5]),
  .I0(sp_inst_0_dout[5]),
  .I1(sp_inst_2_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(dout[6]),
  .I0(sp_inst_0_dout[6]),
  .I1(sp_inst_2_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_23 (
  .O(dout[7]),
  .I0(sp_inst_0_dout[7]),
  .I1(sp_inst_2_dout[7]),
  .S0(dff_q_0)
);
MUX2 mux_inst_26 (
  .O(dout[8]),
  .I0(sp_inst_1_dout[8]),
  .I1(sp_inst_2_dout[8]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(dout[9]),
  .I0(sp_inst_1_dout[9]),
  .I1(sp_inst_2_dout[9]),
  .S0(dff_q_0)
);
MUX2 mux_inst_32 (
  .O(dout[10]),
  .I0(sp_inst_1_dout[10]),
  .I1(sp_inst_2_dout[10]),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(dout[11]),
  .I0(sp_inst_1_dout[11]),
  .I1(sp_inst_2_dout[11]),
  .S0(dff_q_0)
);
MUX2 mux_inst_38 (
  .O(dout[12]),
  .I0(sp_inst_1_dout[12]),
  .I1(sp_inst_2_dout[12]),
  .S0(dff_q_0)
);
MUX2 mux_inst_41 (
  .O(dout[13]),
  .I0(sp_inst_1_dout[13]),
  .I1(sp_inst_2_dout[13]),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(dout[14]),
  .I0(sp_inst_1_dout[14]),
  .I1(sp_inst_2_dout[14]),
  .S0(dff_q_0)
);
MUX2 mux_inst_47 (
  .O(dout[15]),
  .I0(sp_inst_1_dout[15]),
  .I1(sp_inst_2_dout[15]),
  .S0(dff_q_0)
);
MUX2 mux_inst_50 (
  .O(dout[16]),
  .I0(sp_inst_3_dout[16]),
  .I1(sp_inst_5_dout[16]),
  .S0(dff_q_0)
);
MUX2 mux_inst_53 (
  .O(dout[17]),
  .I0(sp_inst_3_dout[17]),
  .I1(sp_inst_5_dout[17]),
  .S0(dff_q_0)
);
MUX2 mux_inst_56 (
  .O(dout[18]),
  .I0(sp_inst_3_dout[18]),
  .I1(sp_inst_5_dout[18]),
  .S0(dff_q_0)
);
MUX2 mux_inst_59 (
  .O(dout[19]),
  .I0(sp_inst_3_dout[19]),
  .I1(sp_inst_5_dout[19]),
  .S0(dff_q_0)
);
MUX2 mux_inst_62 (
  .O(dout[20]),
  .I0(sp_inst_3_dout[20]),
  .I1(sp_inst_5_dout[20]),
  .S0(dff_q_0)
);
MUX2 mux_inst_65 (
  .O(dout[21]),
  .I0(sp_inst_3_dout[21]),
  .I1(sp_inst_5_dout[21]),
  .S0(dff_q_0)
);
MUX2 mux_inst_68 (
  .O(dout[22]),
  .I0(sp_inst_3_dout[22]),
  .I1(sp_inst_5_dout[22]),
  .S0(dff_q_0)
);
MUX2 mux_inst_71 (
  .O(dout[23]),
  .I0(sp_inst_3_dout[23]),
  .I1(sp_inst_5_dout[23]),
  .S0(dff_q_0)
);
MUX2 mux_inst_74 (
  .O(dout[24]),
  .I0(sp_inst_4_dout[24]),
  .I1(sp_inst_5_dout[24]),
  .S0(dff_q_0)
);
MUX2 mux_inst_77 (
  .O(dout[25]),
  .I0(sp_inst_4_dout[25]),
  .I1(sp_inst_5_dout[25]),
  .S0(dff_q_0)
);
MUX2 mux_inst_80 (
  .O(dout[26]),
  .I0(sp_inst_4_dout[26]),
  .I1(sp_inst_5_dout[26]),
  .S0(dff_q_0)
);
MUX2 mux_inst_83 (
  .O(dout[27]),
  .I0(sp_inst_4_dout[27]),
  .I1(sp_inst_5_dout[27]),
  .S0(dff_q_0)
);
MUX2 mux_inst_86 (
  .O(dout[28]),
  .I0(sp_inst_4_dout[28]),
  .I1(sp_inst_5_dout[28]),
  .S0(dff_q_0)
);
MUX2 mux_inst_89 (
  .O(dout[29]),
  .I0(sp_inst_4_dout[29]),
  .I1(sp_inst_5_dout[29]),
  .S0(dff_q_0)
);
MUX2 mux_inst_92 (
  .O(dout[30]),
  .I0(sp_inst_4_dout[30]),
  .I1(sp_inst_5_dout[30]),
  .S0(dff_q_0)
);
MUX2 mux_inst_95 (
  .O(dout[31]),
  .I0(sp_inst_4_dout[31]),
  .I1(sp_inst_5_dout[31]),
  .S0(dff_q_0)
);
endmodule //Gowin_SP_Instr
