module in_dma (
    input clk,
    input rstn,

    input mode_a,
    input mode_b,

    input 
)