`timescale 1ns / 1ps

`include"config.v"
`define USE_INTERNAL_OSC              /*external oscilator not working yet*/
//choose one of USE_CPU_SYSTEM and TEST_DDR
`define USE_CPU_SYSTEM
//`define TEST_DDR
`define TEST_DDR_WITH_AXI_CROSSBAR      /* valid only if TEST_DDR defined. Must choose corresponding GAO manually*/

module TOP # (
    parameter CLK_FREQ = 20_000_000
)(
    input           sys_clk,    //50M
    input           sys_resetn,

    output  [3:0]   led,

    input           RsRx,
    output          RsTx,


    inout   [31:0]  ddr_dq,
    inout   [3:0]   ddr_dqs,
    inout   [3:0]   ddr_dqs_n,
    output  [14:0]  ddr_addr,
    output  [2:0]   ddr_bank,
    output          ddr_cs,
    output          ddr_ras,
    output          ddr_cas,
    output          ddr_we,
    output          ddr_ck,
    output          ddr_ck_n,
    output          ddr_cke,
    output          ddr_odt,
    output          ddr_reset_n,
    output  [3:0]   ddr_dm

    // input            sd_miso,
    // output           sd_clk,
    // output           sd_cs,
    // output           sd_mosi
);

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// clock tree: independent on any reset signals
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

    wire cpu_clk;   /* synthesis syn_keep=1 */ 
    wire core_clk;  /* synthesis syn_keep=1 */ 
    wire ddr_intf_clk;  /* synthesis syn_keep=1 */ 
    wire model_loader_clk;  /* synthesis syn_keep=1 */ 
    wire locked;

    wire ddr_ctl_clk = core_clk;    //use core clk as ddr ctr clock
    wire ddr_ui_clk; /* synthesis syn_keep=1 */ //generated by DDR interface IP core

`ifdef USE_INTERNAL_OSC
    wire clk_osc;   /* synthesis syn_keep=1 */  // 70MHz
    Gowin_OSC OSC_CLOCK(
        .oscout(clk_osc)
    );

    wire clk_20M;   /* synthesis syn_keep=1 */ 
    CLOCK_GEN clk_gen (
        .clk_osc(clk_osc),

        .clk_20M(clk_20M),
        .cpu_clk(cpu_clk),
        .core_clk(core_clk),
        .mem_clk(ddr_intf_clk),
        .model_loader_clk(model_loader_clk),

        .locked(locked)
    );
`else
    Gowin_PLL_ext clk_gen(
        .lock(locked), //output lock
        .clkout0(cpu_clk), // 8M
        .clkout1(ddr_intf_clk), // 200M
        .clkin(sys_clk) //external input 50M
    );
    assign core_clk = sys_clk;
    assign model_loader_clk = sys_clk;
`endif

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// reset tree: sys_resetn input pin triggers all other reset signals
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

    //filter jitter of input sys_resetn
    localparam SYS_RESETN_HIGH_COUNT_MIN = 20'd49999;
    reg [19:0] sys_resetn_counter;
    reg sys_resetn_filtered;/* synthesis syn_keep=1 */
    always @(posedge core_clk or negedge locked) begin
        if (~locked) begin
            sys_resetn_counter <= 0;
            sys_resetn_filtered <= 0;
        end
        else if (~sys_resetn) begin
            sys_resetn_counter <= 0;
            sys_resetn_filtered <= 0;
        end
        else begin
            if (sys_resetn_counter != {20{1'b1}}) begin
                sys_resetn_counter <= sys_resetn_counter + 1'b1;
            end
            sys_resetn_filtered <= sys_resetn_counter >= SYS_RESETN_HIGH_COUNT_MIN;
        end
    end

    //reset sequence for ddr_ui_clk domain
    wire ddr_ui_resetn;     /* synthesis syn_keep=1 */  //generated by DDR controller

    //reset sequence for core_clk domain, triggered by sys_resetn
    wire core_resetn; /* synthesis syn_keep=1 */
    RESET_GEN #(16) core_rst_gen (
        .clk(core_clk),
        .sys_resetn(sys_resetn_filtered),

        .bus_resetn(core_resetn)
    );

    //reset sequence for cpu_clk domain, triggered by sys_resetn
    wire cpu_bus_resetn; /* synthesis syn_keep=1 */
    wire cpu_peri_resetn;/* synthesis syn_keep=1 */
    wire cpu_cpu_resetn; /* synthesis syn_keep=1 */
    RESET_GEN #(16) cpu_rst_gen (
        .clk(cpu_clk),
        .sys_resetn(sys_resetn_filtered),

        .bus_resetn(cpu_bus_resetn),
        .peri_resetn(cpu_peri_resetn),
        .cpu_resetn(cpu_cpu_resetn)
    );

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// network of the main components
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

    wire [31:0]                 fetch_pc;
    wire                        sleeping_o;
    wire                        can_high_freq;
    wire [31:0]                 debug_pc;
    wire [5:0]                  interrupt;

    wire [`CPU_ID_WIDTH  -1 :0] cpu_awid;
    wire [`ADDR_WIDTH    -1 :0] cpu_awaddr;
    wire [`LEN_WIDTH     -1 :0] cpu_awlen;
    wire [`SIZE_WIDTH    -1 :0] cpu_awsize;
    wire [`BURST_WIDTH   -1 :0] cpu_awburst;
    wire [`LOCK_WIDTH    -1 :0] cpu_awlock;
    wire [`CACHE_WIDTH   -1 :0] cpu_awcache;
    wire [`PROT_WIDTH    -1 :0] cpu_awprot;
    wire                        cpu_awvalid;
    wire                        cpu_awready;
    wire [`CPU_ID_WIDTH  -1 :0] cpu_wid;
    wire [`CPU_DATA_WIDTH-1 :0] cpu_wdata;
    wire [`CPU_STRB_WIDTH-1 :0] cpu_wstrb;
    wire                        cpu_wlast;
    wire                        cpu_wvalid;
    wire                        cpu_wready;
    wire [`CPU_ID_WIDTH  -1 :0] cpu_bid;
    wire [`RESP_WIDTH   -1 :0 ] cpu_bresp;
    wire                        cpu_bvalid;
    wire                        cpu_bready;
    wire [`CPU_ID_WIDTH  -1 :0] cpu_arid;
    wire [`ADDR_WIDTH    -1 :0] cpu_araddr;
    wire [`LEN_WIDTH     -1 :0] cpu_arlen;
    wire [`SIZE_WIDTH    -1 :0] cpu_arsize;
    wire [`BURST_WIDTH   -1 :0] cpu_arburst;
    wire [`LOCK_WIDTH    -1 :0] cpu_arlock;
    wire [`CACHE_WIDTH   -1 :0] cpu_arcache;
    wire [`PROT_WIDTH    -1 :0] cpu_arprot;
    wire                        cpu_arvalid;
    wire                        cpu_arready;
    wire [`CPU_ID_WIDTH  -1 :0] cpu_rid;
    wire [`CPU_DATA_WIDTH-1 :0] cpu_rdata;
    wire [`RESP_WIDTH    -1 :0] cpu_rresp;
    wire                        cpu_rlast;
    wire                        cpu_rvalid;
    wire                        cpu_rready;

    wire                        inst_sram_en;
    wire [ 3:0]                 inst_sram_strb;
    wire [31:0]                 inst_sram_wdata;
    wire [31:0]                 inst_sram_rdata;
    wire                        inst_sram_wr;
    wire                        inst_sram_fetch;
    wire [31:0]                 inst_sram_addr;
    wire                        inst_sram_rrdy = 1'b1;
    wire                        inst_sram_ack  = 1'b1;
    wire                        inst_sram_resp = 1'b0;

    wire                        data_sram_en;
    wire [ 3:0]                 data_sram_strb;
    wire [31:0]                 data_sram_wdata;
    wire [31:0]                 data_sram_rdata;
    wire                        data_sram_wr;
    wire                        data_sram_fetch;
    wire [31:0]                 data_sram_addr;
    wire                        data_sram_rrdy = 1'b1;
    wire                        data_sram_ack  = 1'b1;
    wire                        data_sram_resp = 1'b0;

    wire                        timer_int;
    wire                        i2c_int;
    wire                        uart1_int;
    wire                        uart0_int;
    wire                        flash_int;
    wire                        spi_int;
    wire                        vpwm_int;
    wire                        dma_int;

    wire [`ID_WIDTH       -1:0] axi2apb_awid;
    wire [`ADDR_WIDTH    -1 :0] axi2apb_awaddr;
    wire [`LEN_WIDTH     -1 :0] axi2apb_awlen;
    wire [`SIZE_WIDTH    -1 :0] axi2apb_awsize;
    wire [`BURST_WIDTH   -1 :0] axi2apb_awburst;
    wire [`LOCK_WIDTH    -1 :0] axi2apb_awlock;
    wire [`CACHE_WIDTH   -1 :0] axi2apb_awcache;
    wire [`PROT_WIDTH    -1 :0] axi2apb_awprot;
    wire                        axi2apb_awvalid;
    wire                        axi2apb_awready;
    wire [`APB_DATA_WIDTH-1 :0] axi2apb_wdata;
    wire [`APB_STRB_WIDTH-1 :0] axi2apb_wstrb;
    wire                        axi2apb_wlast;
    wire                        axi2apb_wvalid;
    wire                        axi2apb_wready;
    wire [`ID_WIDTH       -1:0] axi2apb_bid;
    wire [`RESP_WIDTH    -1 :0] axi2apb_bresp;
    wire                        axi2apb_bvalid;
    wire                        axi2apb_bready;
    wire [`ID_WIDTH       -1:0] axi2apb_arid;
    wire [`ADDR_WIDTH    -1 :0] axi2apb_araddr;
    wire [`LEN_WIDTH     -1 :0] axi2apb_arlen;
    wire [`SIZE_WIDTH    -1 :0] axi2apb_arsize;
    wire [`BURST_WIDTH   -1 :0] axi2apb_arburst;
    wire [`LOCK_WIDTH    -1 :0] axi2apb_arlock;
    wire [`CACHE_WIDTH   -1 :0] axi2apb_arcache;
    wire [`PROT_WIDTH    -1 :0] axi2apb_arprot;
    wire                        axi2apb_arvalid;
    wire                        axi2apb_arready;
    wire [`ID_WIDTH       -1:0] axi2apb_rid;
    wire [`APB_DATA_WIDTH-1 :0] axi2apb_rdata;
    wire [`RESP_WIDTH    -1 :0] axi2apb_rresp;
    wire                        axi2apb_rlast;
    wire                        axi2apb_rvalid;
    wire                        axi2apb_rready;

    wire                        apb_clk;
    wire                        apb_reset_n;
    wire                        apb_psel;
    wire                        apb_rw;
    wire [`ADDR_WIDTH    -1 :0] apb_addr;
    wire                        apb_enable;
    wire [`APB_DATA_WIDTH-1 :0] apb_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb_datao;
    wire                        apb_ready;

    wire                        apb0_psel;
    wire                        apb0_rw;
    wire [`ADDR_WIDTH    -1 :0] apb0_addr;
    wire                        apb0_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb0_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb0_datao;
    wire                        apb0_ack;

    wire                        apb1_psel;
    wire                        apb1_rw;
    wire [`ADDR_WIDTH    -1 :0] apb1_addr;
    wire                        apb1_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb1_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb1_datao;
    wire                        apb1_ack;

    wire                        apb2_psel;
    wire                        apb2_rw;
    wire [`ADDR_WIDTH    -1 :0] apb2_addr;
    wire                        apb2_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb2_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb2_datao;
    wire                        apb2_ack;

    wire                        apb3_psel;
    wire                        apb3_rw;
    wire [`ADDR_WIDTH    -1 :0] apb3_addr;
    wire                        apb3_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb3_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb3_datao;
    wire                        apb3_ack;

    wire                        apb4_psel;
    wire                        apb4_rw;
    wire [`ADDR_WIDTH    -1 :0] apb4_addr;
    wire                        apb4_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb4_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb4_datao;
    wire                        apb4_ack;

    wire                        apb5_psel;
    wire                        apb5_rw;
    wire [`ADDR_WIDTH    -1 :0] apb5_addr;
    wire                        apb5_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb5_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb5_datao;
    wire                        apb5_ack;

    wire                        apb6_psel;
    wire                        apb6_rw;
    wire [`ADDR_WIDTH    -1 :0] apb6_addr;
    wire                        apb6_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb6_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb6_datao;
    wire                        apb6_ack;

    wire                        apb7_psel;
    wire                        apb7_rw;
    wire [`ADDR_WIDTH    -1 :0] apb7_addr;
    wire                        apb7_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb7_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb7_datao;
    wire                        apb7_ack;

    wire                        apb8_psel;
    wire                        apb8_rw;
    wire [`ADDR_WIDTH    -1 :0] apb8_addr;
    wire                        apb8_enab;
    wire [`APB_DATA_WIDTH-1 :0] apb8_datai;
    wire [`APB_DATA_WIDTH-1 :0] apb8_datao;
    wire                        apb8_ack;

    wire [`ID_WIDTH       -1:0] cpu_ddr_32_awid;
    wire [`ADDR_WIDTH    -1 :0] cpu_ddr_32_awaddr;
    wire [`LEN_WIDTH     -1 :0] cpu_ddr_32_awlen;
    wire [`SIZE_WIDTH    -1 :0] cpu_ddr_32_awsize;
    wire [`BURST_WIDTH   -1 :0] cpu_ddr_32_awburst;
    wire [`LOCK_WIDTH    -1 :0] cpu_ddr_32_awlock;
    wire [`CACHE_WIDTH   -1 :0] cpu_ddr_32_awcache;
    wire [`PROT_WIDTH    -1 :0] cpu_ddr_32_awprot;
    wire                        cpu_ddr_32_awvalid;
    wire                        cpu_ddr_32_awready;
    wire [`DATA_WIDTH    -1 :0] cpu_ddr_32_wdata;
    wire [`STRB_WIDTH    -1 :0] cpu_ddr_32_wstrb;
    wire                        cpu_ddr_32_wlast;
    wire                        cpu_ddr_32_wvalid;
    wire                        cpu_ddr_32_wready;
    wire [`ID_WIDTH       -1:0] cpu_ddr_32_bid;
    wire [`RESP_WIDTH    -1 :0] cpu_ddr_32_bresp;
    wire                        cpu_ddr_32_bvalid;
    wire                        cpu_ddr_32_bready;
    wire [`ID_WIDTH       -1:0] cpu_ddr_32_arid;
    wire [`ADDR_WIDTH    -1 :0] cpu_ddr_32_araddr;
    wire [`LEN_WIDTH     -1 :0] cpu_ddr_32_arlen;
    wire [`SIZE_WIDTH    -1 :0] cpu_ddr_32_arsize;
    wire [`BURST_WIDTH   -1 :0] cpu_ddr_32_arburst;
    wire [`LOCK_WIDTH    -1 :0] cpu_ddr_32_arlock;
    wire [`CACHE_WIDTH   -1 :0] cpu_ddr_32_arcache;
    wire [`PROT_WIDTH    -1 :0] cpu_ddr_32_arprot;
    wire                        cpu_ddr_32_arvalid;
    wire                        cpu_ddr_32_arready;
    wire [`ID_WIDTH       -1:0] cpu_ddr_32_rid;
    wire [`DATA_WIDTH    -1 :0] cpu_ddr_32_rdata;
    wire [`RESP_WIDTH    -1 :0] cpu_ddr_32_rresp;
    wire                        cpu_ddr_32_rlast;
    wire                        cpu_ddr_32_rvalid;
    wire                        cpu_ddr_32_rready;

    wire [`ID_WIDTH       -1:0] cpu_ddr_256_awid;
    wire [`ADDR_WIDTH    -1 :0] cpu_ddr_256_awaddr;
    wire [`LEN_WIDTH     -1 :0] cpu_ddr_256_awlen;
    wire [`SIZE_WIDTH    -1 :0] cpu_ddr_256_awsize;
    wire [`BURST_WIDTH   -1 :0] cpu_ddr_256_awburst;
    wire [`LOCK_WIDTH    -1 :0] cpu_ddr_256_awlock;
    wire [`CACHE_WIDTH   -1 :0] cpu_ddr_256_awcache;
    wire [`PROT_WIDTH    -1 :0] cpu_ddr_256_awprot;
    wire                        cpu_ddr_256_awvalid;
    wire                        cpu_ddr_256_awready;
    wire [`DDR_DATA_WIDTH-1 :0] cpu_ddr_256_wdata;
    wire [`DDR_STRB_WIDTH-1 :0] cpu_ddr_256_wstrb;
    wire                        cpu_ddr_256_wlast;
    wire                        cpu_ddr_256_wvalid;
    wire                        cpu_ddr_256_wready;
    wire [`ID_WIDTH       -1:0] cpu_ddr_256_bid;
    wire [`RESP_WIDTH    -1 :0] cpu_ddr_256_bresp;
    wire                        cpu_ddr_256_bvalid;
    wire                        cpu_ddr_256_bready;
    wire [`ID_WIDTH       -1:0] cpu_ddr_256_arid;
    wire [`ADDR_WIDTH    -1 :0] cpu_ddr_256_araddr;
    wire [`LEN_WIDTH     -1 :0] cpu_ddr_256_arlen;
    wire [`SIZE_WIDTH    -1 :0] cpu_ddr_256_arsize;
    wire [`BURST_WIDTH   -1 :0] cpu_ddr_256_arburst;
    wire [`LOCK_WIDTH    -1 :0] cpu_ddr_256_arlock;
    wire [`CACHE_WIDTH   -1 :0] cpu_ddr_256_arcache;
    wire [`PROT_WIDTH    -1 :0] cpu_ddr_256_arprot;
    wire                        cpu_ddr_256_arvalid;
    wire                        cpu_ddr_256_arready;
    wire [`ID_WIDTH       -1:0] cpu_ddr_256_rid;
    wire [`DDR_DATA_WIDTH-1 :0] cpu_ddr_256_rdata;
    wire [`RESP_WIDTH    -1 :0] cpu_ddr_256_rresp;
    wire                        cpu_ddr_256_rlast;
    wire                        cpu_ddr_256_rvalid;
    wire                        cpu_ddr_256_rready;

    wire [`ID_WIDTH       -1:0] ddr_test_256_awid;
    wire [`ADDR_WIDTH    -1 :0] ddr_test_256_awaddr;
    wire [`LEN_WIDTH     -1 :0] ddr_test_256_awlen;
    wire [`SIZE_WIDTH    -1 :0] ddr_test_256_awsize;
    wire [`BURST_WIDTH   -1 :0] ddr_test_256_awburst;
    wire [`LOCK_WIDTH    -1 :0] ddr_test_256_awlock;
    wire [`CACHE_WIDTH   -1 :0] ddr_test_256_awcache;
    wire [`PROT_WIDTH    -1 :0] ddr_test_256_awprot;
    wire                        ddr_test_256_awvalid;
    wire                        ddr_test_256_awready;
    wire [`DDR_DATA_WIDTH-1 :0] ddr_test_256_wdata;
    wire [`DDR_STRB_WIDTH-1 :0] ddr_test_256_wstrb;
    wire                        ddr_test_256_wlast;
    wire                        ddr_test_256_wvalid;
    wire                        ddr_test_256_wready;
    wire [`ID_WIDTH       -1:0] ddr_test_256_bid;
    wire [`RESP_WIDTH    -1 :0] ddr_test_256_bresp;
    wire                        ddr_test_256_bvalid;
    wire                        ddr_test_256_bready;
    wire [`ID_WIDTH       -1:0] ddr_test_256_arid;
    wire [`ADDR_WIDTH    -1 :0] ddr_test_256_araddr;
    wire [`LEN_WIDTH     -1 :0] ddr_test_256_arlen;
    wire [`SIZE_WIDTH    -1 :0] ddr_test_256_arsize;
    wire [`BURST_WIDTH   -1 :0] ddr_test_256_arburst;
    wire [`LOCK_WIDTH    -1 :0] ddr_test_256_arlock;
    wire [`CACHE_WIDTH   -1 :0] ddr_test_256_arcache;
    wire [`PROT_WIDTH    -1 :0] ddr_test_256_arprot;
    wire                        ddr_test_256_arvalid;
    wire                        ddr_test_256_arready;
    wire [`ID_WIDTH       -1:0] ddr_test_256_rid;
    wire [`DDR_DATA_WIDTH-1 :0] ddr_test_256_rdata;
    wire [`RESP_WIDTH    -1 :0] ddr_test_256_rresp;
    wire                        ddr_test_256_rlast;
    wire                        ddr_test_256_rvalid;
    wire                        ddr_test_256_rready;

    wire [`ID_WIDTH       -1:0] ddr_arb_awid;
    wire [`ADDR_WIDTH    -1 :0] ddr_arb_awaddr;
    wire [7:0]                  ddr_arb_awlen;
    wire [2:0]                  ddr_arb_awsize;
    wire [1:0]                  ddr_arb_awburst;
    wire [1:0]                  ddr_arb_awlock;
    wire [3:0]                  ddr_arb_awcache;
    wire [2:0]                  ddr_arb_awprot;
    wire                        ddr_arb_awvalid;
    wire                        ddr_arb_awready;
    wire [`DDR_DATA_WIDTH-1 :0] ddr_arb_wdata;
    wire [`DDR_STRB_WIDTH-1 :0] ddr_arb_wstrb;
    wire                        ddr_arb_wlast;
    wire                        ddr_arb_wvalid;
    wire                        ddr_arb_wready;
    wire [`ID_WIDTH       -1:0] ddr_arb_bid;
    wire [1:0]                  ddr_arb_bresp;
    wire                        ddr_arb_bvalid;
    wire                        ddr_arb_bready;
    wire [`ID_WIDTH       -1:0] ddr_arb_arid;
    wire [`ADDR_WIDTH    -1 :0] ddr_arb_araddr;
    wire [7:0]                  ddr_arb_arlen;
    wire [2:0]                  ddr_arb_arsize;
    wire [1:0]                  ddr_arb_arburst;
    wire [1:0]                  ddr_arb_arlock;
    wire [3:0]                  ddr_arb_arcache;
    wire [2:0]                  ddr_arb_arprot;
    wire                        ddr_arb_arvalid;
    wire                        ddr_arb_arready;
    wire [`ID_WIDTH       -1:0] ddr_arb_rid;
    wire [`DDR_DATA_WIDTH-1 :0] ddr_arb_rdata;
    wire [1:0]                  ddr_arb_rresp;
    wire                        ddr_arb_rlast;
    wire                        ddr_arb_rvalid;
    wire                        ddr_arb_rready;

    wire                        init_calib_complete;


    wire                        ml_app_rdy;
    wire                        ml_app_cmd_en;
    wire [`ADDR_WIDTH    -1 :0] ml_app_addr;
    wire                        ml_app_wdf_rdy;
    wire [`DATA_WIDTH    -1 :0] ml_app_wdf_data;
    wire [`STRB_WIDTH    -1 :0] ml_app_wdf_mask;
    wire                        ml_app_wdf_wren;

    wire                        init_model_complete;

`ifdef USE_CPU_SYSTEM

    la132_top CPU (
        .boot_pc            (32'h1c000000           ),
        .clk                (cpu_clk                ),
        .clk_count          (cpu_clk                ),
        .hard_resetn        (cpu_cpu_resetn         ),
        .soft_resetn        (cpu_cpu_resetn         ),

        .sleeping           (sleeping_o             ),
        .can_high_freq      (can_high_freq          ),
        .cpu_fetch_pc       (fetch_pc               ),
        .wb_pc              (debug_pc               ),
        .mode_lisa          (1'b1                   ), 
        .inst_xor           (32'b0                  ),

        .nmi                (1'b0                   ),
        .ext_int            (interrupt              ),

        .arid               (cpu_arid[3:0]          ),
        .araddr             (cpu_araddr             ),
        .arlen              (cpu_arlen[3:0]         ),
        .arsize             (cpu_arsize             ),
        .arburst            (cpu_arburst            ),
        .arlock             (cpu_arlock             ),
        .arcache            (cpu_arcache            ),
        .arprot             (cpu_arprot             ),
        .arvalid            (cpu_arvalid            ),
        .arready            (cpu_arready            ),

        .rid                (cpu_rid[3:0]           ),
        .rdata              (cpu_rdata              ),
        .rresp              (cpu_rresp              ),
        .rlast              (cpu_rlast              ),
        .rvalid             (cpu_rvalid             ),
        .rready             (cpu_rready             ),

        .awid               (cpu_awid[3:0]          ),
        .awaddr             (cpu_awaddr             ),
        .awlen              (cpu_awlen[3:0]         ),
        .awsize             (cpu_awsize             ),
        .awburst            (cpu_awburst            ),
        .awlock             (cpu_awlock             ),
        .awcache            (cpu_awcache            ),
        .awprot             (cpu_awprot             ),
        .awvalid            (cpu_awvalid            ),
        .awready            (cpu_awready            ),

        .wid                (cpu_wid[3:0]           ),
        .wdata              (cpu_wdata              ),
        .wstrb              (cpu_wstrb              ),
        .wlast              (cpu_wlast              ),
        .wvalid             (cpu_wvalid             ),
        .wready             (cpu_wready             ),

        .bid                (cpu_bid[3:0]           ),
        .bresp              (cpu_bresp              ),
        .bvalid             (cpu_bvalid             ),
        .bready             (cpu_bready             ),

        .inst_sram_en       (inst_sram_en           ),
        .inst_sram_wr       (inst_sram_wr           ),
        .inst_sram_fetch    (inst_sram_fetch        ),
        .inst_sram_strb     (inst_sram_strb         ),
        .inst_sram_addr     (inst_sram_addr         ),
        .inst_sram_wdata    (inst_sram_wdata        ),
        .inst_sram_rdata    (inst_sram_rdata        ),
        .inst_sram_ack      (inst_sram_ack          ),
        .inst_sram_rrdy     (inst_sram_rrdy         ),
        .inst_sram_resp     (inst_sram_resp         ),

        .data_sram_en       (data_sram_en           ),
        .data_sram_wr       (data_sram_wr           ),
        .data_sram_fetch    (data_sram_fetch        ),
        .data_sram_strb     (data_sram_strb         ),
        .data_sram_addr     (data_sram_addr         ),
        .data_sram_wdata    (data_sram_wdata        ),
        .data_sram_rdata    (data_sram_rdata        ),
        .data_sram_ack      (data_sram_ack          ),
        .data_sram_rrdy     (data_sram_rrdy         ),
        .data_sram_resp     (data_sram_resp         ),

        .trstn              (ljtag_trst_i           ),
        .tck                (ljtag_tck_i            ),
        .tdi                (ljtag_tdi_i            ),
        .tms                (ljtag_tms_i            ),
        .tdo                (ljtag_tdo_o            ),
        .ljtag_prrst        (ljtag_prrst_src        ),
        .ljtag_lock         (1'b0                   ),

        .prid_revision      (4'd0                   ),
        .cpunum             (10'b0                  ),

        .ibus0_valid        (1'b1                   ),
        .ibus0_base         (32'h1c00_0000          ), // va: 1c00_0000 & bfc0_0000
        .ibus0_mask         (32'h1f00_0000          ), // flash 128K, + 4 special page
        .ibus1_valid        (1'b1                   ),
        .ibus1_base         (32'h9f00_0000          ), // va: 9fR0_0000 & bf00_0000
        .ibus1_mask         (32'hdff0_0000          ),
        .ibus2_valid        (1'b0                   ), // flash_en
        .ibus2_base         (32'h9fe6_0000          ), // va: 9fe6_0000 & bfe6_0000
        .ibus2_mask         (32'hdfff_ff00          ),
        .ibus3_valid        (1'b0                   ), // compact_mem&flash_en),
        .ibus3_base         (32'h8000_3000          ), // for va: 8000_30xx & 0000_00xx -> pa: 0000_30xx & 4000_00xx
        .ibus3_mask         (32'h7fff_ff00          ),
        .dbus0_valid        (1'b1                   ),
        .dbus0_base         (32'h8000_0000          ),
        .dbus0_mask         (32'hdfff_e000          ), // 8K byte, for va: 8000_0000 & a000_0000 -> pa: 0000_0000
        .dbus1_valid        (1'b1                   ),
        .dbus1_base         (32'h0000_0000          ),
        .dbus1_mask         (32'hffff_e000          ), // 8K byte, for va: 0000_0000             -> pa: 0000_0000
        .dbus2_valid        (1'b0                   ), // unused
        .dbus2_base         (32'h0000_0000          ),
        .dbus2_mask         (32'h0000_0000          ),
        .dbus3_valid        (1'b0                   ), // unused
        .dbus3_base         (32'h0000_0000          ),
        .dbus3_mask         (32'h0000_0000          ),

        .test_mode          (1'b0                   )
    );

    Gowin_SP_Instr IRAM (
        .dout               (inst_sram_rdata        ), //output [31:0] dout
        .clk                (cpu_clk                ), //input clk
        .oce                (inst_sram_en           ), //input oce
        .ce                 (inst_sram_en           ), //input ce
        .reset              (~cpu_peri_resetn       ), //input reset
        .wre                (inst_sram_wr           ), //input wre
        .ad                 (inst_sram_addr[13:2]   ), //input [11:0] ad
        .din                (inst_sram_wdata        ) //input [31:0] din
    );


    Gowin_SP_Data DRAM (
        .dout               (data_sram_rdata        ), //output [31:0] dout
        .clk                (cpu_clk                ), //input clk
        .oce                (data_sram_en           ), //input oce
        .ce                 (data_sram_en           ), //input ce
        .reset              (~cpu_peri_resetn       ), //input reset
        .wre                (data_sram_wr           ), //input wre
        .ad                 (data_sram_addr[13:2]   ), //input [11:0] ad
        .din                (data_sram_wdata        ) //input [31:0] din
    );

    axicb_crossbar_top # (
        .AXI_ADDR_W         (`ADDR_WIDTH            ),
        .AXI_ID_W           (`ID_WIDTH              ),
        .AXI_DATA_W         (`DATA_WIDTH            ),
        .AXI_SIGNALING      (1                      ),
        .USER_SUPPORT       (1                      ),

        .MST0_CDC           (1                      ),
        .MST0_ID_MASK       ('h20                   ),
        .MST0_OSTDREQ_NUM   (0                      ),
        .MST0_PRIORITY      (0                      ),

        .SLV0_CDC           (0                      ),
        .SLV0_START_ADDR    (`APB_ADDR_BASE         ),
        .SLV0_END_ADDR      (`APB_ADDR_END          ),
        .SLV0_OSTDREQ_NUM   (0                      ),
        .SLV0_KEEP_BASE_ADDR(1                      ),

        .SLV1_CDC           (0                      ),
        .SLV1_START_ADDR    (`DDR_ADDR_BASE         ),
        .SLV1_END_ADDR      (`DDR_ADDR_END          ),
        .SLV1_OSTDREQ_NUM   (0                      ),
        .SLV1_KEEP_BASE_ADDR(1                      )
    ) AXI_crossbar_32 (
        .aclk               (core_clk               ),
        .aresetn            (core_resetn            ),
        .srst               (~core_resetn           ),
        .slv0_aclk          (cpu_clk                ),
        .slv0_aresetn       (cpu_bus_resetn         ),
        .slv0_srst          (~cpu_bus_resetn        ),////////////////////////////
        .slv0_awvalid       (cpu_awvalid            ),
        .slv0_awready       (cpu_awready            ),
        .slv0_awaddr        (cpu_awaddr             ),
        .slv0_awlen         (cpu_awlen              ),
        .slv0_awsize        (cpu_awsize             ),
        .slv0_awburst       (cpu_awburst            ),
        .slv0_awlock        (cpu_awlock             ),
        .slv0_awcache       (cpu_awcache            ),
        .slv0_awprot        (cpu_awprot             ),
        .slv0_awid          ({4'h2,cpu_awid}        ),
        .slv0_wvalid        (cpu_wvalid             ),
        .slv0_wready        (cpu_wready             ),
        .slv0_wlast         (cpu_wlast              ),
        .slv0_wdata         (cpu_wdata              ),
        .slv0_wstrb         (cpu_wstrb              ),
        .slv0_bvalid        (cpu_bvalid             ),
        .slv0_bready        (cpu_bready             ),
        .slv0_bid           (cpu_bid                ),
        .slv0_bresp         (cpu_bresp              ),
        .slv0_arvalid       (cpu_arvalid            ),
        .slv0_arready       (cpu_arready            ),
        .slv0_araddr        (cpu_araddr             ),
        .slv0_arlen         (cpu_arlen              ),
        .slv0_arsize        (cpu_arsize             ),
        .slv0_arburst       (cpu_arburst            ),
        .slv0_arlock        (cpu_arlock             ),
        .slv0_arcache       (cpu_arcache            ),
        .slv0_arprot        (cpu_arprot             ),
        .slv0_arid          ({4'h2,cpu_arid}        ),
        .slv0_rvalid        (cpu_rvalid             ),
        .slv0_rready        (cpu_rready             ),
        .slv0_rid           (cpu_rid                ),
        .slv0_rresp         (cpu_rresp              ),
        .slv0_rdata         (cpu_rdata              ),
        .slv0_rlast         (cpu_rlast              ),

        .mst0_aclk          (core_clk               ),
        .mst0_aresetn       (core_resetn            ),
        .mst0_srst          (~core_resetn           ),
        .mst0_awvalid       (axi2apb_awvalid        ),
        .mst0_awready       (axi2apb_awready        ),
        .mst0_awaddr        (axi2apb_awaddr         ),
        .mst0_awlen         (axi2apb_awlen          ),
        .mst0_awsize        (axi2apb_awsize         ),
        .mst0_awburst       (axi2apb_awburst        ),
        .mst0_awlock        (axi2apb_awlock         ),
        .mst0_awcache       (axi2apb_awcache        ),
        .mst0_awprot        (axi2apb_awprot         ),
        .mst0_awid          (axi2apb_awid           ),
        .mst0_wvalid        (axi2apb_wvalid         ),
        .mst0_wready        (axi2apb_wready         ),
        .mst0_wlast         (axi2apb_wlast          ),
        .mst0_wdata         (axi2apb_wdata          ),
        .mst0_wstrb         (axi2apb_wstrb          ),
        .mst0_bvalid        (axi2apb_bvalid         ),
        .mst0_bready        (axi2apb_bready         ),
        .mst0_bid           (axi2apb_bid            ),
        .mst0_bresp         (axi2apb_bresp          ),
        .mst0_arvalid       (axi2apb_arvalid        ),
        .mst0_arready       (axi2apb_arready        ),
        .mst0_araddr        (axi2apb_araddr         ),
        .mst0_arlen         (axi2apb_arlen          ),
        .mst0_arsize        (axi2apb_arsize         ),
        .mst0_arburst       (axi2apb_arburst        ),
        .mst0_arlock        (axi2apb_arlock         ),
        .mst0_arcache       (axi2apb_arcache        ),
        .mst0_arprot        (axi2apb_arprot         ),
        .mst0_arid          (axi2apb_arid           ),
        .mst0_rvalid        (axi2apb_rvalid         ),
        .mst0_rready        (axi2apb_rready         ),
        .mst0_rid           (axi2apb_rid            ),
        .mst0_rresp         (axi2apb_rresp          ),
        .mst0_rdata         (axi2apb_rdata          ),
        .mst0_rlast         (axi2apb_rlast          ),

        .mst1_aclk          (core_clk               ),
        .mst1_aresetn       (core_resetn            ),
        .mst1_srst          (~core_resetn           ),
        .mst1_awvalid       (cpu_ddr_32_awvalid        ),
        .mst1_awready       (cpu_ddr_32_awready        ),
        .mst1_awaddr        (cpu_ddr_32_awaddr         ),
        .mst1_awlen         (cpu_ddr_32_awlen          ),
        .mst1_awsize        (cpu_ddr_32_awsize         ),
        .mst1_awburst       (cpu_ddr_32_awburst        ),
        .mst1_awlock        (cpu_ddr_32_awlock         ),
        .mst1_awcache       (cpu_ddr_32_awcache        ),
        .mst1_awprot        (cpu_ddr_32_awprot         ),
        .mst1_awid          (cpu_ddr_32_awid           ),
        .mst1_wvalid        (cpu_ddr_32_wvalid         ),
        .mst1_wready        (cpu_ddr_32_wready         ),
        .mst1_wlast         (cpu_ddr_32_wlast          ),
        .mst1_wdata         (cpu_ddr_32_wdata          ),
        .mst1_wstrb         (cpu_ddr_32_wstrb          ),
        .mst1_bvalid        (cpu_ddr_32_bvalid         ),
        .mst1_bready        (cpu_ddr_32_bready         ),
        .mst1_bid           (cpu_ddr_32_bid            ),
        .mst1_bresp         (cpu_ddr_32_bresp          ),
        .mst1_arvalid       (cpu_ddr_32_arvalid        ),
        .mst1_arready       (cpu_ddr_32_arready        ),
        .mst1_araddr        (cpu_ddr_32_araddr         ),
        .mst1_arlen         (cpu_ddr_32_arlen          ),
        .mst1_arsize        (cpu_ddr_32_arsize         ),
        .mst1_arburst       (cpu_ddr_32_arburst        ),
        .mst1_arlock        (cpu_ddr_32_arlock         ),
        .mst1_arcache       (cpu_ddr_32_arcache        ),
        .mst1_arprot        (cpu_ddr_32_arprot         ),
        .mst1_arid          (cpu_ddr_32_arid           ),
        .mst1_rvalid        (cpu_ddr_32_rvalid         ),
        .mst1_rready        (cpu_ddr_32_rready         ),
        .mst1_rid           (cpu_ddr_32_rid            ),
        .mst1_rresp         (cpu_ddr_32_rresp          ),
        .mst1_rdata         (cpu_ddr_32_rdata          ),
        .mst1_rlast         (cpu_ddr_32_rlast          )
    );

    axi_adapter # (
        .ADDR_WIDTH         (`ADDR_WIDTH            ),
        .S_DATA_WIDTH       (`DATA_WIDTH            ),
        .M_DATA_WIDTH       (`DDR_DATA_WIDTH        )
    ) axi_adapter_32_to_256 (
        .clk                (core_clk               ),
        .rst                (~core_resetn           ),

        .s_axi_awid         (cpu_ddr_32_awid        ),
        .s_axi_awaddr       (cpu_ddr_32_awaddr      ),
        .s_axi_awlen        (cpu_ddr_32_awlen       ),
        .s_axi_awsize       (cpu_ddr_32_awsize      ),
        .s_axi_awburst      (cpu_ddr_32_awburst     ),
        .s_axi_awlock       (cpu_ddr_32_awlock      ),
        .s_axi_awcache      (cpu_ddr_32_awcache     ),
        .s_axi_awprot       (cpu_ddr_32_awprot      ),
        .s_axi_awvalid      (cpu_ddr_32_awvalid     ),
        .s_axi_awready      (cpu_ddr_32_awready     ),
        .s_axi_wdata        (cpu_ddr_32_wdata       ),
        .s_axi_wstrb        (cpu_ddr_32_wstrb       ),
        .s_axi_wlast        (cpu_ddr_32_wlast       ),
        .s_axi_wvalid       (cpu_ddr_32_wvalid      ),
        .s_axi_wready       (cpu_ddr_32_wready      ),
        .s_axi_bid          (cpu_ddr_32_bid         ),
        .s_axi_bresp        (cpu_ddr_32_bresp       ),
        .s_axi_bvalid       (cpu_ddr_32_bvalid      ),
        .s_axi_bready       (cpu_ddr_32_bready      ),
        .s_axi_arid         (cpu_ddr_32_arid        ),
        .s_axi_araddr       (cpu_ddr_32_araddr      ),
        .s_axi_arlen        (cpu_ddr_32_arlen       ),
        .s_axi_arsize       (cpu_ddr_32_arsize      ),
        .s_axi_arburst      (cpu_ddr_32_arburst     ),
        .s_axi_arlock       (cpu_ddr_32_arlock      ),
        .s_axi_arcache      (cpu_ddr_32_arcache     ),
        .s_axi_arprot       (cpu_ddr_32_arprot      ),
        .s_axi_arvalid      (cpu_ddr_32_arvalid     ),
        .s_axi_arready      (cpu_ddr_32_arready     ),
        .s_axi_rid          (cpu_ddr_32_rid         ),
        .s_axi_rdata        (cpu_ddr_32_rdata       ),
        .s_axi_rresp        (cpu_ddr_32_rresp       ),
        .s_axi_rlast        (cpu_ddr_32_rlast       ),
        .s_axi_rvalid       (cpu_ddr_32_rvalid      ),
        .s_axi_rready       (cpu_ddr_32_rready      ),
    
        .m_axi_awid         (cpu_ddr_256_awid       ),
        .m_axi_awaddr       (cpu_ddr_256_awaddr     ),
        .m_axi_awlen        (cpu_ddr_256_awlen      ),
        .m_axi_awsize       (cpu_ddr_256_awsize     ),
        .m_axi_awburst      (cpu_ddr_256_awburst    ),
        .m_axi_awlock       (cpu_ddr_256_awlock     ),
        .m_axi_awcache      (cpu_ddr_256_awcache    ),
        .m_axi_awprot       (cpu_ddr_256_awprot     ),
        .m_axi_awvalid      (cpu_ddr_256_awvalid    ),
        .m_axi_awready      (cpu_ddr_256_awready    ),
        .m_axi_wdata        (cpu_ddr_256_wdata      ),
        .m_axi_wstrb        (cpu_ddr_256_wstrb      ),
        .m_axi_wlast        (cpu_ddr_256_wlast      ),
        .m_axi_wvalid       (cpu_ddr_256_wvalid     ),
        .m_axi_wready       (cpu_ddr_256_wready     ),
        .m_axi_bid          (cpu_ddr_256_bid        ),
        .m_axi_bresp        (cpu_ddr_256_bresp      ),
        .m_axi_bvalid       (cpu_ddr_256_bvalid     ),
        .m_axi_bready       (cpu_ddr_256_bready     ),
        .m_axi_arid         (cpu_ddr_256_arid       ),
        .m_axi_araddr       (cpu_ddr_256_araddr     ),
        .m_axi_arlen        (cpu_ddr_256_arlen      ),
        .m_axi_arsize       (cpu_ddr_256_arsize     ),
        .m_axi_arburst      (cpu_ddr_256_arburst    ),
        .m_axi_arlock       (cpu_ddr_256_arlock     ),
        .m_axi_arcache      (cpu_ddr_256_arcache    ),
        .m_axi_arprot       (cpu_ddr_256_arprot     ),
        .m_axi_arvalid      (cpu_ddr_256_arvalid    ),
        .m_axi_arready      (cpu_ddr_256_arready    ),
        .m_axi_rid          (cpu_ddr_256_rid        ),
        .m_axi_rdata        (cpu_ddr_256_rdata      ),
        .m_axi_rresp        (cpu_ddr_256_rresp      ),
        .m_axi_rlast        (cpu_ddr_256_rlast      ),
        .m_axi_rvalid       (cpu_ddr_256_rvalid     ),
        .m_axi_rready       (cpu_ddr_256_rready     )
    );

    /*
     * AXI-32 SLAVE 0
     */
    axi2apb_bridge #(
        .ID_WIDTH           (`ID_WIDTH              ),
        .ADDR_WIDTH         (`ADDR_WIDTH            ),
        .DATA_WIDTH         (`APB_DATA_WIDTH        )
    ) apb (
        .clk                (core_clk               ),
        .rst_n              (core_resetn            ),
        .axi_s_awid         (axi2apb_awid           ),
        .axi_s_awaddr       (axi2apb_awaddr         ),
        .axi_s_awlen        (axi2apb_awlen          ),
        .axi_s_awsize       (axi2apb_awsize         ),
        .axi_s_awburst      (axi2apb_awburst        ),
        .axi_s_awlock       (axi2apb_awlock         ),
        .axi_s_awcache      (axi2apb_awcache        ),
        .axi_s_awprot       (axi2apb_awprot         ),
        .axi_s_awvalid      (axi2apb_awvalid        ),
        .axi_s_awready      (axi2apb_awready        ),

        .axi_s_wid          (axi2apb_awid           ),
        .axi_s_wdata        (axi2apb_wdata          ),
        .axi_s_wstrb        (axi2apb_wstrb          ),
        .axi_s_wlast        (axi2apb_wlast          ),
        .axi_s_wvalid       (axi2apb_wvalid         ),
        .axi_s_wready       (axi2apb_wready         ),

        .axi_s_bid          (axi2apb_bid            ),
        .axi_s_bresp        (axi2apb_bresp          ),
        .axi_s_bvalid       (axi2apb_bvalid         ),
        .axi_s_bready       (axi2apb_bready         ),

        .axi_s_arid         (axi2apb_arid           ),
        .axi_s_araddr       (axi2apb_araddr         ),
        .axi_s_arlen        (axi2apb_arlen          ),
        .axi_s_arsize       (axi2apb_arsize         ),
        .axi_s_arburst      (axi2apb_arburst        ),
        .axi_s_arlock       (axi2apb_arlock         ),
        .axi_s_arcache      (axi2apb_arcache        ),
        .axi_s_arprot       (axi2apb_arprot         ),
        .axi_s_arvalid      (axi2apb_arvalid        ),
        .axi_s_arready      (axi2apb_arready        ),

        .axi_s_rid          (axi2apb_rid            ),
        .axi_s_rdata        (axi2apb_rdata          ),
        .axi_s_rresp        (axi2apb_rresp          ),
        .axi_s_rlast        (axi2apb_rlast          ),
        .axi_s_rvalid       (axi2apb_rvalid         ),
        .axi_s_rready       (axi2apb_rready         ),

        .apb_clk            (apb_clk                ),
        .apb_reset_n        (apb_reset_n            ),
        .reg_psel           (apb_psel               ),
        .reg_rw             (apb_rw                 ),
        .reg_addr           (apb_addr               ),
        .reg_enable         (apb_enable             ),
        .reg_datai          (apb_datai              ),
        .reg_datao          (apb_datao              ),
        .reg_ready_1        (apb_ready              )
    );


    apb_mux9 apb_mux (
        .apb_psel_cpu       (apb_psel               ),
        .apb_rw_cpu         (apb_rw                 ),
        .apb_addr_cpu       (apb_addr               ),
        .apb_enab_cpu       (apb_enable             ),
        .apb_datai_cpu      (apb_datai              ),
        .apb_datao_cpu      (apb_datao              ),
        .apb_ack_cpu        (apb_ready              ),

        .apb0_psel          (apb0_psel              ),
        .apb0_rw            (apb0_rw                ),
        .apb0_addr          (apb0_addr              ),
        .apb0_enab          (apb0_enab              ),
        .apb0_datai         (apb0_datai             ),
        .apb0_datao         (apb0_datao             ),
        .apb0_ack           (apb0_ack               ),

        .apb1_psel          (apb1_psel              ),
        .apb1_rw            (apb1_rw                ),
        .apb1_addr          (apb1_addr              ),
        .apb1_enab          (apb1_enab              ),
        .apb1_datai         (apb1_datai             ),
        .apb1_datao         (apb1_datao             ),
        .apb1_ack           (apb1_ack               ),
        
        .apb2_psel          (apb2_psel              ),
        .apb2_rw            (apb2_rw                ),
        .apb2_addr          (apb2_addr              ),
        .apb2_enab          (apb2_enab              ),
        .apb2_datai         (apb2_datai             ),
        .apb2_datao         (apb2_datao             ),
        .apb2_ack           (apb2_ack               ),
        
        .apb3_psel          (apb3_psel              ),
        .apb3_rw            (apb3_rw                ),
        .apb3_addr          (apb3_addr              ),
        .apb3_enab          (apb3_enab              ),
        .apb3_datai         (apb3_datai             ),
        .apb3_datao         (apb3_datao             ),
        .apb3_ack           (apb3_ack               ),
        
        .apb4_psel          (apb4_psel              ),
        .apb4_rw            (apb4_rw                ),
        .apb4_addr          (apb4_addr              ),
        .apb4_enab          (apb4_enab              ),
        .apb4_datai         (apb4_datai             ),
        .apb4_datao         (apb4_datao             ),
        .apb4_ack           (apb4_ack               ),
        
        .apb5_psel          (apb5_psel              ),
        .apb5_rw            (apb5_rw                ),
        .apb5_addr          (apb5_addr              ),
        .apb5_enab          (apb5_enab              ),
        .apb5_datai         (apb5_datai             ),
        .apb5_datao         (apb5_datao             ),
        .apb5_ack           (apb5_ack               ),
        
        .apb6_psel          (apb6_psel              ),
        .apb6_rw            (apb6_rw                ),
        .apb6_addr          (apb6_addr              ),
        .apb6_enab          (apb6_enab              ),
        .apb6_datai         (apb6_datai             ),
        .apb6_datao         (apb6_datao             ),
        .apb6_ack           (apb6_ack               ),
        
        .apb7_psel          (apb7_psel              ),
        .apb7_rw            (apb7_rw                ),
        .apb7_addr          (apb7_addr              ),
        .apb7_enab          (apb7_enab              ),
        .apb7_datai         (apb7_datai             ),
        .apb7_datao         (apb7_datao             ),
        .apb7_ack           (apb7_ack               ),
        
        .apb8_psel          (apb8_psel              ),
        .apb8_rw            (apb8_rw                ),
        .apb8_addr          (apb8_addr              ),
        .apb8_enab          (apb8_enab              ),
        .apb8_datai         (apb8_datai             ),
        .apb8_datao         (apb8_datao             ),
        .apb8_ack           (apb8_ack               )
    );
    
    CONFREG IntController(
        .apb_pclk           (apb_clk                ),
        .apb_prstn          (apb_reset_n            ),
        
        .apb_psel           (apb0_psel              ),
        .apb_pwrite         (apb0_rw                ),
        .apb_paddr          (apb0_addr              ),
        .apb_penable        (apb0_enab              ),
        .apb_pwdata         (apb0_datai             ),
        .apb_prdata         (apb0_datao             ),
        .apb_ack            (apb0_ack               ),

        .timer_int          (timer_int              ),
        .i2c_int            (i2c_int                ),
        .uart1_int          (uart1_int              ),
        .uart0_int          (uart0_int              ),
        .flash_int          (flash_int              ),
        .spi_int            (spi_int                ),
        .vpwm_int           (vpwm_int               ),
        .dma_int            (dma_int                ),

        .int_o              (interrupt[4]           )
    );
    
    UART_TOP # (
        .CLK_FREQ           (50_000_000             )
    ) UART1 (
        .apb_pclk           (apb_clk                ),
        .apb_prstn          (apb_reset_n            ),

        .apb_psel           (apb1_psel              ),
        .apb_pwrite         (apb1_rw                ),
        .apb_paddr          (apb1_addr              ),
        .apb_penable        (apb1_enab              ),
        .apb_pwdata         (apb1_datai             ),
        .apb_prdata         (apb1_datao             ),
        .uart_ready         (apb1_ack               ),

        .RsRx               (RsRx                   ),
        .RsTx               (RsTx                   ),
        .uart_irq           (uart1_int              )
    );

    
    LED_driver LED (
        .clk                (apb_clk                ),
        .resetn             (apb_reset_n            ),
        .apb_psel           (apb8_psel              ),
        .apb_rw             (apb8_rw                ),
        .apb_addr           (apb8_addr              ),
        .apb_enab           (apb8_enab              ),
        .apb_datai          (apb8_datai             ),
        .apb_datao          (apb8_datao             ),
        .apb_ack            (apb8_ack               ),

        .led                (led[3:1]               )
    );

`endif

`ifdef TEST_DDR
`ifdef TEST_DDR_WITH_AXI_CROSSBAR
    ddr_ctr_wr_rd_test test(
        .clk                (core_clk                   ),//crossing into ddr_ui_clk by AXI crossbar
        .rstn               (core_resetn                ),
        
        .awaddr             (ddr_test_256_awaddr         ),
        .awid               (ddr_test_256_awid           ),
        .awvalid            (ddr_test_256_awvalid        ),
        .awburst            (ddr_test_256_awburst        ),
        .awsize             (ddr_test_256_awsize         ),
        .awlen              (ddr_test_256_awlen          ),
        .awready            (ddr_test_256_awready        ),
        .wdata              (ddr_test_256_wdata          ),
        .wstrb              (ddr_test_256_wstrb          ),
        .wlast              (ddr_test_256_wlast          ),
        .wvalid             (ddr_test_256_wvalid         ),
        .wready             (ddr_test_256_wready         ),
        .bvalid             (ddr_test_256_bvalid         ),
        .bready             (ddr_test_256_bready         ),
        .araddr             (ddr_test_256_araddr         ),
        .arid               (ddr_test_256_arid           ),
        .arvalid            (ddr_test_256_arvalid        ),
        .arburst            (ddr_test_256_arburst        ),
        .arsize             (ddr_test_256_arsize         ),
        .arlen              (ddr_test_256_arlen          ),
        .arready            (ddr_test_256_arready        ),
        .rdata              (ddr_test_256_rdata          ),
        .rvalid             (ddr_test_256_rvalid         ),
        .rready             (ddr_test_256_rready         ),

        .led                (led[1]                 ),

        .ddr_ready          (init_calib_complete    )
    );

`else
    ddr_ctr_wr_rd_test test(
        .clk                (ddr_ui_clk             ),//directly attached to ddr_ui_clk
        .rstn               (ddr_ui_resetn          ),
        
        .awaddr             (ddr_arb_awaddr         ),
        .awid               (ddr_arb_awid           ),
        .awvalid            (ddr_arb_awvalid        ),
        .awburst            (ddr_arb_awburst        ),
        .awsize             (ddr_arb_awsize         ),
        .awlen              (ddr_arb_awlen          ),
        .awready            (ddr_arb_awready        ),
        .wdata              (ddr_arb_wdata          ),
        .wstrb              (ddr_arb_wstrb          ),
        .wlast              (ddr_arb_wlast          ),
        .wvalid             (ddr_arb_wvalid         ),
        .wready             (ddr_arb_wready         ),
        .bvalid             (ddr_arb_bvalid         ),
        .bready             (ddr_arb_bready         ),
        .araddr             (ddr_arb_araddr         ),
        .arid               (ddr_arb_arid           ),
        .arvalid            (ddr_arb_arvalid        ),
        .arburst            (ddr_arb_arburst        ),
        .arsize             (ddr_arb_arsize         ),
        .arlen              (ddr_arb_arlen          ),
        .arready            (ddr_arb_arready        ),
        .rdata              (ddr_arb_rdata          ),
        .rvalid             (ddr_arb_rvalid         ),
        .rready             (ddr_arb_rready         ),

        .led                (led[1]                 ),

        .ddr_ready          (init_calib_complete    )
     );

`endif
`endif

`ifndef TEST_DDR
`define USE_AXI_256_CROSSBAR
`else
`ifdef TEST_DDR_WITH_AXI_CROSSBAR
`define USE_AXI_256_CROSSBAR
`endif
`endif

`ifdef USE_AXI_256_CROSSBAR
    axicb_crossbar_top # (
        .AXI_ADDR_W         (`ADDR_WIDTH            ),
        .AXI_ID_W           (`ID_WIDTH      ),
        .AXI_DATA_W         (`DDR_DATA_WIDTH        ),

        .AXI_SIGNALING      (1                      ),
        .USER_SUPPORT       (1                      ),

        .MST0_CDC           (0                      ),
        .MST0_ID_MASK       ('h10                   ),
        .MST0_OSTDREQ_NUM   (0                      ),
        .MST0_PRIORITY      (0                      ),

        .MST1_CDC           (0                      ),
        .MST1_ID_MASK       ('h20                   ),
        .MST1_OSTDREQ_NUM   (0                      ),
        .MST1_PRIORITY      (0                      ),
        
        .MST2_CDC           (0                      ),
        .MST2_ID_MASK       ('h40                   ),
        .MST2_OSTDREQ_NUM   (0                      ),
        .MST2_PRIORITY      (0                      ),

        .SLV0_CDC           (1                      ),
        .SLV0_START_ADDR    (`DDR_ADDR_BASE         ),
        .SLV0_END_ADDR      (`DDR_ADDR_END          ),
        .SLV0_OSTDREQ_NUM   (0                      ),
        .SLV0_KEEP_BASE_ADDR(1                      )
    ) AXI_crossbar_256 (
        .aclk               (core_clk               ),
        .aresetn            (1'b1                   ),
        .srst               (~core_resetn           ),

        .slv0_aclk          (core_clk               ),
        .slv0_aresetn       (1'b1                   ),
        .slv0_srst          (~core_resetn           ),////////////////////////////
        .slv0_awvalid       (ddr_test_256_awvalid   ),
        .slv0_awready       (ddr_test_256_awready   ),
        .slv0_awaddr        (ddr_test_256_awaddr    ),
        .slv0_awlen         (ddr_test_256_awlen     ),
        .slv0_awsize        (ddr_test_256_awsize    ),
        .slv0_awburst       (ddr_test_256_awburst   ),
        .slv0_awlock        (ddr_test_256_awlock    ),
        .slv0_awcache       (ddr_test_256_awcache   ),
        .slv0_awprot        (ddr_test_256_awprot    ),
        .slv0_awid          (ddr_test_256_awid      ),
        .slv0_wvalid        (ddr_test_256_wvalid    ),
        .slv0_wready        (ddr_test_256_wready    ),
        .slv0_wlast         (ddr_test_256_wlast     ),
        .slv0_wdata         (ddr_test_256_wdata     ),
        .slv0_wstrb         (ddr_test_256_wstrb     ),
        .slv0_bvalid        (ddr_test_256_bvalid    ),
        .slv0_bready        (ddr_test_256_bready    ),
        .slv0_bid           (ddr_test_256_bid       ),
        .slv0_bresp         (ddr_test_256_bresp     ),
        .slv0_arvalid       (ddr_test_256_arvalid   ),
        .slv0_arready       (ddr_test_256_arready   ),
        .slv0_araddr        (ddr_test_256_araddr    ),
        .slv0_arlen         (ddr_test_256_arlen     ),
        .slv0_arsize        (ddr_test_256_arsize    ),
        .slv0_arburst       (ddr_test_256_arburst   ),
        .slv0_arlock        (ddr_test_256_arlock    ),
        .slv0_arcache       (ddr_test_256_arcache   ),
        .slv0_arprot        (ddr_test_256_arprot    ),
        .slv0_arid          (ddr_test_256_arid      ),
        .slv0_rvalid        (ddr_test_256_rvalid    ),
        .slv0_rready        (ddr_test_256_rready    ),
        .slv0_rid           (ddr_test_256_rid       ),
        .slv0_rresp         (ddr_test_256_rresp     ),
        .slv0_rdata         (ddr_test_256_rdata     ),
        .slv0_rlast         (ddr_test_256_rlast     ),

        .slv1_aclk          (core_clk               ),
        .slv1_aresetn       (1'b1                   ),
        .slv1_srst          (~core_resetn           ),////////////////////////////
        .slv1_awvalid       (cpu_ddr_256_awvalid    ),
        .slv1_awready       (cpu_ddr_256_awready    ),
        .slv1_awaddr        (cpu_ddr_256_awaddr     ),
        .slv1_awlen         (cpu_ddr_256_awlen      ),
        .slv1_awsize        (cpu_ddr_256_awsize     ),
        .slv1_awburst       (cpu_ddr_256_awburst    ),
        .slv1_awlock        (cpu_ddr_256_awlock     ),
        .slv1_awcache       (cpu_ddr_256_awcache    ),
        .slv1_awprot        (cpu_ddr_256_awprot     ),
        .slv1_awid          (cpu_ddr_256_awid       ),
        .slv1_wvalid        (cpu_ddr_256_wvalid     ),
        .slv1_wready        (cpu_ddr_256_wready     ),
        .slv1_wlast         (cpu_ddr_256_wlast      ),
        .slv1_wdata         (cpu_ddr_256_wdata      ),
        .slv1_wstrb         (cpu_ddr_256_wstrb      ),
        .slv1_bvalid        (cpu_ddr_256_bvalid     ),
        .slv1_bready        (cpu_ddr_256_bready     ),
        .slv1_bid           (cpu_ddr_256_bid        ),
        .slv1_bresp         (cpu_ddr_256_bresp      ),
        .slv1_arvalid       (cpu_ddr_256_arvalid    ),
        .slv1_arready       (cpu_ddr_256_arready    ),
        .slv1_araddr        (cpu_ddr_256_araddr     ),
        .slv1_arlen         (cpu_ddr_256_arlen      ),
        .slv1_arsize        (cpu_ddr_256_arsize     ),
        .slv1_arburst       (cpu_ddr_256_arburst    ),
        .slv1_arlock        (cpu_ddr_256_arlock     ),
        .slv1_arcache       (cpu_ddr_256_arcache    ),
        .slv1_arprot        (cpu_ddr_256_arprot     ),
        .slv1_arid          (cpu_ddr_256_arid       ),
        .slv1_rvalid        (cpu_ddr_256_rvalid     ),
        .slv1_rready        (cpu_ddr_256_rready     ),
        .slv1_rid           (cpu_ddr_256_rid        ),
        .slv1_rresp         (cpu_ddr_256_rresp      ),
        .slv1_rdata         (cpu_ddr_256_rdata      ),
        .slv1_rlast         (cpu_ddr_256_rlast      ),

        .mst0_aclk          (ddr_ui_clk             ),
        .mst0_aresetn       (1'b1                   ),
        .mst0_srst          (~ddr_ui_resetn         ),
        .mst0_awvalid       (ddr_arb_awvalid        ),
        .mst0_awready       (ddr_arb_awready        ),
        .mst0_awaddr        (ddr_arb_awaddr         ),
        .mst0_awlen         (ddr_arb_awlen          ),
        .mst0_awsize        (ddr_arb_awsize         ),
        .mst0_awburst       (ddr_arb_awburst        ),
        .mst0_awlock        (ddr_arb_awlock         ),
        .mst0_awcache       (ddr_arb_awcache        ),
        .mst0_awprot        (ddr_arb_awprot         ),
        .mst0_awid          (ddr_arb_awid           ),
        .mst0_wvalid        (ddr_arb_wvalid         ),
        .mst0_wready        (ddr_arb_wready         ),
        .mst0_wlast         (ddr_arb_wlast          ),
        .mst0_wdata         (ddr_arb_wdata          ),
        .mst0_wstrb         (ddr_arb_wstrb          ),
        .mst0_bvalid        (ddr_arb_bvalid         ),
        .mst0_bready        (ddr_arb_bready         ),
        .mst0_bid           (ddr_arb_bid            ),
        .mst0_bresp         (ddr_arb_bresp          ),
        .mst0_arvalid       (ddr_arb_arvalid        ),
        .mst0_arready       (ddr_arb_arready        ),
        .mst0_araddr        (ddr_arb_araddr         ),
        .mst0_arlen         (ddr_arb_arlen          ),
        .mst0_arsize        (ddr_arb_arsize         ),
        .mst0_arburst       (ddr_arb_arburst        ),
        .mst0_arlock        (ddr_arb_arlock         ),
        .mst0_arcache       (ddr_arb_arcache        ),
        .mst0_arprot        (ddr_arb_arprot         ),
        .mst0_arid          (ddr_arb_arid           ),
        .mst0_rvalid        (ddr_arb_rvalid         ),
        .mst0_rready        (ddr_arb_rready         ),
        .mst0_rid           (ddr_arb_rid            ),
        .mst0_rresp         (ddr_arb_rresp          ),
        .mst0_rdata         (ddr_arb_rdata          ),
        .mst0_rlast         (ddr_arb_rlast          )
    );
`endif

    /*
     * AXI-256 SLAVE 0
     */
    DDR_Controller # (
        .DATA_WIDTH         (`DDR_DATA_WIDTH        ),
        .ADDR_WIDTH         (`ADDR_WIDTH            ),
        .ID_WIDTH           (`ID_WIDTH              ),
        .AXI_ID             (8'h10                  )
    ) ddr_ctr (
        .ctr_clk            (ddr_ctl_clk            ),
        .memory_clk         (ddr_intf_clk           ),
        .pll_lock           (locked                 ),
        .sys_resetn         (sys_resetn_filtered    ),
        .axi_aresetn        (ddr_ui_resetn          ),
        .ui_clk             (ddr_ui_clk             ),
        .ui_sync_resetn     (ddr_ui_resetn          ),
        .init_calib_complete(init_calib_complete    ),

        .s_axi_awid         (ddr_arb_awid           ),
        .s_axi_awaddr       (ddr_arb_awaddr         ),
        .s_axi_awlen        (ddr_arb_awlen          ),
        .s_axi_awsize       (ddr_arb_awsize         ),
        .s_axi_awburst      (ddr_arb_awburst        ),
        .s_axi_awlock       (ddr_arb_awlock[0]      ),
        .s_axi_awcache      (ddr_arb_awcache        ),
        .s_axi_awprot       (ddr_arb_awprot         ),
        .s_axi_awvalid      (ddr_arb_awvalid        ),
        .s_axi_awready      (ddr_arb_awready        ),
        .s_axi_wdata        (ddr_arb_wdata          ),
        .s_axi_wstrb        (ddr_arb_wstrb          ),
        .s_axi_wlast        (ddr_arb_wlast          ),
        .s_axi_wvalid       (ddr_arb_wvalid         ),
        .s_axi_wready       (ddr_arb_wready         ),
        .s_axi_bid          (ddr_arb_bid            ),
        .s_axi_bresp        (ddr_arb_bresp          ),
        .s_axi_bvalid       (ddr_arb_bvalid         ),
        .s_axi_bready       (ddr_arb_bready         ),
        .s_axi_arid         (ddr_arb_arid           ),
        .s_axi_araddr       (ddr_arb_araddr         ),
        .s_axi_arlen        (ddr_arb_arlen          ),
        .s_axi_arsize       (ddr_arb_arsize         ),
        .s_axi_arburst      (ddr_arb_arburst        ),
        .s_axi_arlock       (ddr_arb_arlock[0]      ),
        .s_axi_arcache      (ddr_arb_arcache        ),
        .s_axi_arprot       (ddr_arb_arprot         ),
        .s_axi_arvalid      (ddr_arb_arvalid        ),
        .s_axi_arready      (ddr_arb_arready        ),
        .s_axi_rid          (ddr_arb_rid            ),
        .s_axi_rdata        (ddr_arb_rdata          ),
        .s_axi_rresp        (ddr_arb_rresp          ),
        .s_axi_rlast        (ddr_arb_rlast          ),
        .s_axi_ruser        (ddr_arb_ruser          ),
        .s_axi_rvalid       (ddr_arb_rvalid         ),
        .s_axi_rready       (ddr_arb_rready         ),

        .ddr_dq             (ddr_dq                 ),
        .ddr_dqs            (ddr_dqs                ),
        .ddr_dqs_n          (ddr_dqs_n              ),
        .ddr_addr           (ddr_addr               ),
        .ddr_bank           (ddr_bank               ),
        .ddr_cs             (ddr_cs                 ),
        .ddr_ras            (ddr_ras                ),
        .ddr_cas            (ddr_cas                ),
        .ddr_we             (ddr_we                 ),
        .ddr_ck             (ddr_ck                 ),
        .ddr_ck_n           (ddr_ck_n               ),
        .ddr_cke            (ddr_cke                ),
        .ddr_odt            (ddr_odt                ),
        .ddr_reset_n        (ddr_reset_n            ),
        .ddr_dm             (ddr_dm                 )
    );
    // assign led[2:0] = 0;
    assign led[0] = ~init_calib_complete;

    assign init_model_complete = 1'b1;

endmodule

