//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.01 (64-bit)
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Thu Mar 28 21:38:10 2024

module Gowin_SP_Instr (dout, clk, oce, ce, reset, wre, ad, din);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [13:0] ad;
input [31:0] din;

wire lut_f_0;
wire [26:0] spx9_inst_0_dout_w;
wire [8:0] spx9_inst_0_dout;
wire [26:0] spx9_inst_1_dout_w;
wire [8:0] spx9_inst_1_dout;
wire [26:0] spx9_inst_2_dout_w;
wire [8:0] spx9_inst_2_dout;
wire [26:0] spx9_inst_3_dout_w;
wire [8:0] spx9_inst_3_dout;
wire [26:0] spx9_inst_4_dout_w;
wire [17:9] spx9_inst_4_dout;
wire [26:0] spx9_inst_5_dout_w;
wire [17:9] spx9_inst_5_dout;
wire [26:0] spx9_inst_6_dout_w;
wire [17:9] spx9_inst_6_dout;
wire [26:0] spx9_inst_7_dout_w;
wire [17:9] spx9_inst_7_dout;
wire [29:0] sp_inst_8_dout_w;
wire [19:18] sp_inst_8_dout;
wire [29:0] sp_inst_9_dout_w;
wire [21:20] sp_inst_9_dout;
wire [29:0] sp_inst_10_dout_w;
wire [23:22] sp_inst_10_dout;
wire [29:0] sp_inst_11_dout_w;
wire [25:24] sp_inst_11_dout;
wire [29:0] sp_inst_12_dout_w;
wire [27:26] sp_inst_12_dout;
wire [29:0] sp_inst_13_dout_w;
wire [29:28] sp_inst_13_dout;
wire [29:0] sp_inst_14_dout_w;
wire [31:30] sp_inst_14_dout;
wire [27:0] sp_inst_15_dout_w;
wire [3:0] sp_inst_15_dout;
wire [27:0] sp_inst_16_dout_w;
wire [7:4] sp_inst_16_dout;
wire [27:0] sp_inst_17_dout_w;
wire [11:8] sp_inst_17_dout;
wire [27:0] sp_inst_18_dout_w;
wire [15:12] sp_inst_18_dout;
wire [27:0] sp_inst_19_dout_w;
wire [19:16] sp_inst_19_dout;
wire [27:0] sp_inst_20_dout_w;
wire [23:20] sp_inst_20_dout;
wire [27:0] sp_inst_21_dout_w;
wire [27:24] sp_inst_21_dout;
wire [27:0] sp_inst_22_dout_w;
wire [31:28] sp_inst_22_dout;
wire [31:0] sp_inst_23_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire mux_o_12;
wire mux_o_13;
wire mux_o_16;
wire mux_o_17;
wire mux_o_31;
wire mux_o_32;
wire mux_o_35;
wire mux_o_36;
wire mux_o_50;
wire mux_o_51;
wire mux_o_54;
wire mux_o_55;
wire mux_o_69;
wire mux_o_70;
wire mux_o_73;
wire mux_o_74;
wire mux_o_88;
wire mux_o_89;
wire mux_o_92;
wire mux_o_93;
wire mux_o_107;
wire mux_o_108;
wire mux_o_111;
wire mux_o_112;
wire mux_o_126;
wire mux_o_127;
wire mux_o_130;
wire mux_o_131;
wire mux_o_145;
wire mux_o_146;
wire mux_o_149;
wire mux_o_150;
wire mux_o_164;
wire mux_o_165;
wire mux_o_168;
wire mux_o_169;
wire mux_o_183;
wire mux_o_184;
wire mux_o_187;
wire mux_o_188;
wire mux_o_202;
wire mux_o_203;
wire mux_o_206;
wire mux_o_207;
wire mux_o_221;
wire mux_o_222;
wire mux_o_225;
wire mux_o_226;
wire mux_o_240;
wire mux_o_241;
wire mux_o_244;
wire mux_o_245;
wire mux_o_259;
wire mux_o_260;
wire mux_o_263;
wire mux_o_264;
wire mux_o_278;
wire mux_o_279;
wire mux_o_282;
wire mux_o_283;
wire mux_o_297;
wire mux_o_298;
wire mux_o_301;
wire mux_o_302;
wire mux_o_316;
wire mux_o_317;
wire mux_o_320;
wire mux_o_321;
wire mux_o_335;
wire mux_o_336;
wire mux_o_339;
wire mux_o_340;
wire mux_o_352;
wire mux_o_364;
wire mux_o_376;
wire mux_o_388;
wire mux_o_400;
wire mux_o_412;
wire mux_o_424;
wire mux_o_436;
wire mux_o_448;
wire mux_o_460;
wire mux_o_472;
wire mux_o_484;
wire mux_o_496;
wire mux_o_508;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

LUT5 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[9]),
  .I1(ad[10]),
  .I2(ad[11]),
  .I3(ad[12]),
  .I4(ad[13])
);
defparam lut_inst_0.INIT = 32'h01000000;
SPX9 spx9_inst_0 (
    .DO({spx9_inst_0_dout_w[26:0],spx9_inst_0_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_0.READ_MODE = 1'b0;
defparam spx9_inst_0.WRITE_MODE = 2'b01;
defparam spx9_inst_0.BIT_WIDTH = 9;
defparam spx9_inst_0.BLK_SEL = 3'b000;
defparam spx9_inst_0.RESET_MODE = "SYNC";
defparam spx9_inst_0.INIT_RAM_00 = 288'hC67B3198C160B0182C166B31980D66B41B8C0673F1DEF17E3059AD07E401FF0F7DBC000D;
defparam spx9_inst_0.INIT_RAM_01 = 288'h0000000000000000000000000000000000000000000001000040003188F000C16630D82C;
defparam spx9_inst_0.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_0.INIT_RAM_20 = 288'hD0637418DD0637418DD063418A350AAD54A95429D4CA5522D166B258AC15EAE56AB0AA35;
defparam spx9_inst_0.INIT_RAM_21 = 288'h52A9168B3592C560AF572B5585500003418D000000000000000000000000000D0637418D;
defparam spx9_inst_0.INIT_RAM_22 = 288'hFF813218CC62B38085078381AC603184C620C20323F0884020001551A8556AA54AA14EA6;
defparam spx9_inst_0.INIT_RAM_23 = 288'h582BD5CAD561546A208FC221008FFCA5D8078FC221008C04B1122031987FE04FFF3BDFAD;
defparam spx9_inst_0.INIT_RAM_24 = 288'hC66B01A00CA85558B65128D42AB552A550A75329548BF5F2F578BB5D2E570B75A2CD64B1;
defparam spx9_inst_0.INIT_RAM_25 = 288'h552A550A75329548BF5F2F578BB5D2E570B75A2CD64B1582BD5CAD56157FE8402003599F;
defparam spx9_inst_0.INIT_RAM_26 = 288'h6660319AC6633400C06663198C06030198C656310EC7631880198C060B16AB65128D42AB;
defparam spx9_inst_0.INIT_RAM_27 = 288'h3B18C40633B0031ACD6663418CD6663198CCD633758CC66B3358CD0633199AC66035998C;
defparam spx9_inst_0.INIT_RAM_28 = 288'hC6EB75BCC663381A006067F198CC603001AC66B31998C666375A0CD6B319A00603158876;
defparam spx9_inst_0.INIT_RAM_29 = 288'h6031588763B18C40633B0031BADD6F319D8C660373F8CC66301800C6B331B8C6633318CC;
defparam spx9_inst_0.INIT_RAM_2A = 288'h066B598CDC6EB75BCC663381B9FC6633180C00001818D06335998C666375A0CD6B319A00;
defparam spx9_inst_0.INIT_RAM_2B = 288'h006B19ACC66631998DD6EB798CC670373F8CC66301800006B19ACC6663198CCC63331BAD;
defparam spx9_inst_0.INIT_RAM_2C = 288'h06637180C3B1D8C620319D8018DD6F341A0CC7630198DD6EB4198DC6030EC7631880C676;
defparam spx9_inst_0.INIT_RAM_2D = 288'h319D8C384667FFFF8402B33FECC06300EC763098C40633B0031BADD68331B8C066375BAD;
defparam spx9_inst_0.INIT_RAM_2E = 288'h3B18401FFFFE100ACCFFFFD980C601D8EC6131880C676308033F8C467FC00763B184C620;
defparam spx9_inst_0.INIT_RAM_2F = 288'h3B1D8C2631018CEC61C263199FFFFE100ACCFFE100ACCFFB0180C066030EC763098C4063;
defparam spx9_inst_0.INIT_RAM_30 = 288'h1018CEC61007FFFFFFC201599FFFFB3318CC6663198CCC6331998C6633318CC6603180C4;
defparam spx9_inst_0.INIT_RAM_31 = 288'h62FFF0805667FFFECCC6331998C6633318CC6663198CCC6331980C603198AC43B1D8C263;
defparam spx9_inst_0.INIT_RAM_32 = 288'h6633318CC6663198CCC6331998C6633018C06331588763B184C620319D8C200FFFFFFEC4;
defparam spx9_inst_0.INIT_RAM_33 = 288'h31880C676308000004C2B31988C3B1D8C2631018CEC61007FFFEC462FFF0805667FD998C;
defparam spx9_inst_0.INIT_RAM_34 = 288'h66EB39ACE66F300F80D73359800603319800FF811980C6660199806631D8CC5621D8EC61;
defparam spx9_inst_0.INIT_RAM_35 = 288'h06335980C0063358CDC63331ACC6680199CCC673B5ACE66B333ECC6663198CC03E8398CE;
defparam spx9_inst_0.INIT_RAM_36 = 288'hD60319A00621D8EC6131880C67630E10180C6633318CCFFE13198CC6330018CC6631998D;
defparam spx9_inst_0.INIT_RAM_37 = 288'h6632D94C96431D8CC5621D8EC6131880C67630E10199F6633318CC6663199FFC2333FE04;
defparam spx9_inst_0.INIT_RAM_38 = 288'hC6333018CD6632598DD6037198CD633718CC66033580C66B3319AC66B3000C066331998C;
defparam spx9_inst_0.INIT_RAM_39 = 288'h6633318CCFFE118A0603E3198006663198CCC6333FF84C663198006663198CCC6333FF84;
defparam spx9_inst_0.INIT_RAM_3A = 288'h66001998C6633318CCFFE118A0603E3198006663198CCC6333FF84628180F8C66001998C;
defparam spx9_inst_0.INIT_RAM_3B = 288'h6663199FF02001998C6633318CCFFE118A0603E3198006663198CCC6333FF84628180F8C;
defparam spx9_inst_0.INIT_RAM_3C = 288'hC6EB19B8C66634198DD633718CC6663198CCD663319CC6763199AD0633400C0666319800;
defparam spx9_inst_0.INIT_RAM_3D = 288'h0663758CDC63331A0CC6EB19B8C6633318CC666B3198CE633B18CCD68319A00607FF1A0C;
defparam spx9_inst_0.INIT_RAM_3E = 288'h621D8EC631018CEC61C20333F8CD633598CCC6333FF84667FC09AC063340000FF813FF8D;
defparam spx9_inst_0.INIT_RAM_3F = 288'h06B3300CCC6B331B8CC66319980666341ACCC6835998D66637580CC6E31998D06B3180C0;

SPX9 spx9_inst_1 (
    .DO({spx9_inst_1_dout_w[26:0],spx9_inst_1_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_1.READ_MODE = 1'b0;
defparam spx9_inst_1.WRITE_MODE = 2'b01;
defparam spx9_inst_1.BIT_WIDTH = 9;
defparam spx9_inst_1.BLK_SEL = 3'b001;
defparam spx9_inst_1.RESET_MODE = "SYNC";
defparam spx9_inst_1.INIT_RAM_00 = 288'hC0030EC7631880C676006359ACCCFE33198C6600198AC621D8EC631018CEC0066631998D;
defparam spx9_inst_1.INIT_RAM_01 = 288'h3B18C40633B000580C3B1D8C620319D800203B1D8C620319D8018C061D8EC631018CEC00;
defparam spx9_inst_1.INIT_RAM_02 = 288'h66E3018CCD6337598CF6637180C6033318CCC033188763B18C40633B00059AC063358876;
defparam spx9_inst_1.INIT_RAM_03 = 288'h00333198CC6031988C3B1D8C620319D8018DE6837180CC76301800C6EB7180CC6E30198D;
defparam spx9_inst_1.INIT_RAM_04 = 288'h6663198CCC6333FF84667FC09AC0633400C43B1D8C2631018CEC00C6B3419AC0663718CC;
defparam spx9_inst_1.INIT_RAM_05 = 288'h66B3000C06633001FF0233018CCC033300CC63B198AC43B1D8C2631018CEC61C20333ECC;
defparam spx9_inst_1.INIT_RAM_06 = 288'h6663598CD00333998CE76B59CCD6667D98CCC63319807D07319CCDD67359CCDE601F01AE;
defparam spx9_inst_1.INIT_RAM_07 = 288'h1018CEC61C203018CC6663199FFC2633198C66003198CC63331A0C66B301800C66B19B8C;
defparam spx9_inst_1.INIT_RAM_08 = 288'h66E3198CC066B018CD6663358CD6600180CC6633318CC65B2992C863B198AC43B1D8C263;
defparam spx9_inst_1.INIT_RAM_09 = 288'hC6331998C667FF098CC633000CCC6331998C667FF098C6660319ACC64331BAC06E3319AC;
defparam spx9_inst_1.INIT_RAM_0A = 288'hC633000CCC6331998C667FF08C50301F18CC0033318CC6663199FFC23140C07C633000CC;
defparam spx9_inst_1.INIT_RAM_0B = 288'hC23140C07C633000CCC6331998C667FF08C50301F18CC0033318CC6663199FFC23140C07;
defparam spx9_inst_1.INIT_RAM_0C = 288'hC633199ACC663398CEC63335A0C6680180CCC633000CCC6333FE040033318CC6663199FF;
defparam spx9_inst_1.INIT_RAM_0D = 288'h6663198CCD663319CC6763199AD0633400C0FFE34198DD633718CCC68331BAC66E3198CC;
defparam spx9_inst_1.INIT_RAM_0E = 288'hE60359D80667FF08CCFF813580C6680001FF027FF1A0CC6EB19B8C66634198DD633718CC;
defparam spx9_inst_1.INIT_RAM_0F = 288'h3B1D8C620319D8C3840667F19AC66B31998C6667D9B8D66000000000001998C566000FA0;
defparam spx9_inst_1.INIT_RAM_10 = 288'h66310EC763098C40633B003180C3B1D8C620319D80180061D8EC631018CED846633018C0;
defparam spx9_inst_1.INIT_RAM_11 = 288'h006B318CCC6B33598C66635998D66237FEC43B1D8C2631018CEC6100635988DFFE019980;
defparam spx9_inst_1.INIT_RAM_12 = 288'h66B13FF8466003FF84667FD80C060310EC763098C40633B18709ACC63335ACDC6331980C;
defparam spx9_inst_1.INIT_RAM_13 = 288'hC26B3182C66B10EC763098C40633B18401FFC263198C43B1D8C2631018CEC61007FF58CC;
defparam spx9_inst_1.INIT_RAM_14 = 288'hC06319B8D660018AC43B1D8C620319D8C200FFE13580C66B10EC763098C40633B18401FF;
defparam spx9_inst_1.INIT_RAM_15 = 288'h66633190C6030188763B18C40633B613598C6633318CCC6E3199ACC633B1CCCC6B30000C;
defparam spx9_inst_1.INIT_RAM_16 = 288'h66635998DC663318CCC6B331B8CC63331ACCC6E33198C66635998DC663318CC66633190C;
defparam spx9_inst_1.INIT_RAM_17 = 288'h666341ACCC0631998D0663598C43B1D8C620319D8018D66637198CC63331ACCC6E33198C;
defparam spx9_inst_1.INIT_RAM_18 = 288'h0663999ADC67B00F80E78331CCCC6F300F80D70331ACCC6836198D06B33018C66634198D;
defparam spx9_inst_1.INIT_RAM_19 = 288'hC663199ADC67B00F80E78331CCCC6E31998DC64331BED03E839E0DD7337598CF601F01CF;
defparam spx9_inst_1.INIT_RAM_1A = 288'h31880C67630803FEC4007FD8980663318A8C3B1D8C2631018CEC00C6837190CC6E3219AD;
defparam spx9_inst_1.INIT_RAM_1B = 288'h006375A0CC7731980EC6830018DD68331C0CE63301D8D0660198CC6663418CD62B10EC76;
defparam spx9_inst_1.INIT_RAM_1C = 288'h3B1D8C620319D8018DD68331DCC6603B1A0C006375A0CC703398CC0763419806633318CC;
defparam spx9_inst_1.INIT_RAM_1D = 288'hC6330018DD68331DCC6603B1A0C006375A0CC703398CC07634198066331998D063358AC4;
defparam spx9_inst_1.INIT_RAM_1E = 288'hC6030EC7631880C676006375A0CC7731980EC6830018DD68331C0CE63301D8D0660198CC;
defparam spx9_inst_1.INIT_RAM_1F = 288'hC60331D8C066379BADF6E30198EC6033018C663018AC43B1D8C620319D8018DD6EB4198D;
defparam spx9_inst_1.INIT_RAM_20 = 288'h66635998D666B718CCC6B331ACCD6E31998D660031ACCD683318CCC6B33018C666379A0D;
defparam spx9_inst_1.INIT_RAM_21 = 288'hC6B335B8C66635998D666B4198C666359800C6B335B8C6663599AC06635998D666B4198C;
defparam spx9_inst_1.INIT_RAM_22 = 288'h31880C67600601998D06B331A0D6660198C43B1D8C620319D8018D666B4198C666359800;
defparam spx9_inst_1.INIT_RAM_23 = 288'h319D8018DE6B34198E063331BAD5683188763B18C40633B0031ACCD6B331ACC62B10EC76;
defparam spx9_inst_1.INIT_RAM_24 = 288'h6601F41CC67635998D06B31998C163018AC43B1D8C2631018CEC00C6EB55A0C3B1D8C620;
defparam spx9_inst_1.INIT_RAM_25 = 288'h6660318CCC6B331BAC06637598C66637598C66635998D6663718CCC6B331ACC6663318CC;
defparam spx9_inst_1.INIT_RAM_26 = 288'hC03331A0D666341ACCC6835998DD6C3598C43B1D8C620319D8C200000131ACCC6B331A0D;
defparam spx9_inst_1.INIT_RAM_27 = 288'h31880C67600635998DD60331B8C660031ACCC6E33198C6660198C5621D8EC631018CEC00;
defparam spx9_inst_1.INIT_RAM_28 = 288'hC63331ACC003118CC5621D8EC6131880C676308031A0D066359ACC0031198AC621D8EC61;
defparam spx9_inst_1.INIT_RAM_29 = 288'h423930ACC6663199806600188CCD63319AAC621D8EC6131880C676308031ACCC6E3319AC;
defparam spx9_inst_1.INIT_RAM_2A = 288'hC633000CCC633188763B18C40633B184018D068331ACD667FD08E4C2B3199AC0633401FF;
defparam spx9_inst_1.INIT_RAM_2B = 288'h3B184C620319D8018D66637198CC6333018C6633318CC621D8EC631018CEC00CFE3198CC;
defparam spx9_inst_1.INIT_RAM_2C = 288'hC663019FF027FC098503333FE84726174CCD66333198CC663198CCC633199AC662B51876;
defparam spx9_inst_1.INIT_RAM_2D = 288'hFF8130ACCFFA11C980C6633180CFF813FE04C2E3199FF423930ACC6663199FF42393018C;
defparam spx9_inst_1.INIT_RAM_2E = 288'hC663198CCC6331988C3B1D8C2631018CEC61007FC09FF02017FE8472603198CC6033FE04;
defparam spx9_inst_1.INIT_RAM_2F = 288'h6633318CCFFA11C985667FD08E4C0633198C067FC09FF026140CCCFFA11C98566333198C;
defparam spx9_inst_1.INIT_RAM_30 = 288'h020140DFF42393018CC663019FF027FC098503333FE8472603198CC6033FE04FF8130B8C;
defparam spx9_inst_1.INIT_RAM_31 = 288'h006B018CD66633180C00333198C066341B8C061D8EC631018CEC61C2331998C067FC09FF;
defparam spx9_inst_1.INIT_RAM_32 = 288'h66E359B8C066379BADF6B3819AC06335998CC603000CCC663018C662B10EC7631880C676;
defparam spx9_inst_1.INIT_RAM_33 = 288'hE6633D98EC63335B8CC63331B8C66310EC7631880C676006341B8C060031A0DC6033580C;
defparam spx9_inst_1.INIT_RAM_34 = 288'hD6F30198EC63331B8C66310EC7631880C67600637188CD6E3318CCD6F33182CC763199AD;
defparam spx9_inst_1.INIT_RAM_35 = 288'hF663B18CCC6E3198C43B1D8C620319D8018DC62331BAD66EB3198CC63335BCC0663B18CC;
defparam spx9_inst_1.INIT_RAM_36 = 288'hC663199ADC663318CCD6E33198C666B7198CC63335B8CC663199ADE63B31D8C666B7998C;
defparam spx9_inst_1.INIT_RAM_37 = 288'h319D8018DE6837180CC76301800C6EB7180CC6E30198066310EC7631880C6760063519AD;
defparam spx9_inst_1.INIT_RAM_38 = 288'hC66B3188CC6E3198CC461D8EC631018CED84C6633198CD6631198DC6331988C3B1D8C620;
defparam spx9_inst_1.INIT_RAM_39 = 288'h31880C676006375A8CC6A30EC7631880C676006375A8CC6A30EC7631880C676C2633198C;
defparam spx9_inst_1.INIT_RAM_3A = 288'h3B18C40633B003598CF6EB51BAFD6B375DAD66E3319ACC62331B8C6633358CC56A30EC76;
defparam spx9_inst_1.INIT_RAM_3B = 288'h3B184C620319D801ACE67B75A8DD7EB59B8CC66B3188CC6E31998EC633199AC662B51876;
defparam spx9_inst_1.INIT_RAM_3C = 288'h66031980C66230EC763098C40633B184018D06335998C667FF09A566E319800603311876;
defparam spx9_inst_1.INIT_RAM_3D = 288'h66031980C6033018CC0633019FFC2331980C66031980C6033019FFC2331980C66031980C;
defparam spx9_inst_1.INIT_RAM_3E = 288'h467FF098C6600180763B184C620319D8C200FF813FF846667F198C46003FFFFC233180C0;
defparam spx9_inst_1.INIT_RAM_3F = 288'hC68319ACCC6333FE847261719AC66E319800607FD08E4C68319ACCC63331BCC67631998D;

SPX9 spx9_inst_2 (
    .DO({spx9_inst_2_dout_w[26:0],spx9_inst_2_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_2.READ_MODE = 1'b0;
defparam spx9_inst_2.WRITE_MODE = 2'b01;
defparam spx9_inst_2.BIT_WIDTH = 9;
defparam spx9_inst_2.BLK_SEL = 3'b010;
defparam spx9_inst_2.RESET_MODE = "SYNC";
defparam spx9_inst_2.INIT_RAM_00 = 288'hC60331BAD66E301980C6033000C621D8EC631018CEC61007FD08E4C2B31998CC6633188C;
defparam spx9_inst_2.INIT_RAM_01 = 288'h06635998E066379A0CC6B331C0CC6EB75A0CC6E301980C63331BCD06635998E066375ACD;
defparam spx9_inst_2.INIT_RAM_02 = 288'h666375A6D666375A2D666341ACCC6835998D06B331BAD16B3188763B18C40633B0031BCD;
defparam spx9_inst_2.INIT_RAM_03 = 288'hC033188763B18C40633B0031BAD066341800C6EB4198D0660198C43B1D8C620319D80180;
defparam spx9_inst_2.INIT_RAM_04 = 288'h3B18C40633B0031BADE6834198EC60331BAD066341800C6EB75A0CC6E30198DD68331A0C;
defparam spx9_inst_2.INIT_RAM_05 = 288'h06637198C066379ACD0663818C43B1D8C620319DB08CC60001980CC06B1998D063018876;
defparam spx9_inst_2.INIT_RAM_06 = 288'h621D8EC631018CEC61000010984C2B331A0DC6631988C3B1D8C2631018CEC00C6EB75B8C;
defparam spx9_inst_2.INIT_RAM_07 = 288'h6663718CCC6B331ACCC6E319980666B318CCC6B331ACCC6E31998D66E335ACDC633198AC;
defparam spx9_inst_2.INIT_RAM_08 = 288'h3B184C620319DB080062B10EC7631880C6760060199ACC63331ACCC6B331B8C66635998D;
defparam spx9_inst_2.INIT_RAM_09 = 288'h66B3318CCFFA11C9C5C3633598C666B59B8E6600181FF4239001AC06337580C66B158876;
defparam spx9_inst_2.INIT_RAM_0A = 288'hC63335ACDC0233FEC4C2E33598C666B59A006033318CC0067D19FF423130B8CD663199AD;
defparam spx9_inst_2.INIT_RAM_0B = 288'h6261719ACC63335ACD666319800FFA11C9C5F361F19ACC63335ACDC7EB318CCD6B371DAC;
defparam spx9_inst_2.INIT_RAM_0C = 288'h31880C67630E101800007FD08C4007FD08C4C0233FE846261719ACC63335ACDCFA33FE84;
defparam spx9_inst_2.INIT_RAM_0D = 288'h66000000000001998C567FD08C4CFB371ACC0000000000033318ECC6837180CFF9D8EC61;
defparam spx9_inst_2.INIT_RAM_0E = 288'h002B51800D2E13198DC63333ECDC6B3000000000000CCC62B3FE8462315998C6667D9B8D;
defparam spx9_inst_2.INIT_RAM_0F = 288'h0033318ACFFA11898566330199F66E3598000000000006663159FF423118ACCC6231988C;
defparam spx9_inst_2.INIT_RAM_10 = 288'hC61B3FE0402E7D9B8D66000000000001998C367FFFE0402FFC0805CFB371ACC000000000;
defparam spx9_inst_2.INIT_RAM_11 = 288'h66E3418CD62B10EC763098C40633B61018763B18FFFFF020173ECDC6B3000000000000CC;
defparam spx9_inst_2.INIT_RAM_12 = 288'h66E0318CC00301988C00613198C66001980CD60319AC400613198C6600019FF423131A0C;
defparam spx9_inst_2.INIT_RAM_13 = 288'h621D8EC6131880C67630E1019AC66335998C667FD08C4C2E3319AC66337FE846261758CC;
defparam spx9_inst_2.INIT_RAM_14 = 288'h603311800C263318CC0033019AC063358800C263318CC00033FE846263418CDC68319AC5;
defparam spx9_inst_2.INIT_RAM_15 = 288'h30E1019AC66335998C667FD08C4C2E3358CCC6E3199FF423130BAC6663718CCC06319800;
defparam spx9_inst_2.INIT_RAM_16 = 288'h66B31988C00613198C663100184C66319800067FD08C4D60319AC5621D8EC6131880C676;
defparam spx9_inst_2.INIT_RAM_17 = 288'h00613198C663100184C66319800067FD08C4D60319AC5621D8EC6131880C67630E10198D;
defparam spx9_inst_2.INIT_RAM_18 = 288'h66033580CC6E3199AC0663718CCD60331ACC60310EC763098C40633B187080CC6B3598C4;
defparam spx9_inst_2.INIT_RAM_19 = 288'h66803580C66EB018CDD60319ACCC66B198CD0033018C00033018CC066B0198D66001980C;
defparam spx9_inst_2.INIT_RAM_1A = 288'h063371A0C66801998CD63335ACC66E3418CDC68319A006663358CCD6B319B8D063371A0C;
defparam spx9_inst_2.INIT_RAM_1B = 288'hFFA1188006663358CCD6B319BAC66E31998D063340000FFA1188006663358CCD6B319B8D;
defparam spx9_inst_2.INIT_RAM_1C = 288'hC66319800067FD08C4D60319AC5621D8EC6131880C67630E11999FC66B198CD666319800;
defparam spx9_inst_2.INIT_RAM_1D = 288'h42310EC763098C40633B187080CFFA1189FF623140DFF42313FEC4FFE13198C66313FF84;
defparam spx9_inst_2.INIT_RAM_1E = 288'hD6631198DC633000C0FFA1189FF423130B8CC6233FE8462617198C467FD08C4C2E3119FF;
defparam spx9_inst_2.INIT_RAM_1F = 288'h42310EC763098C40633B187080CC68319ACCC6333FE84623174D87C6733188CC7631998D;
defparam spx9_inst_2.INIT_RAM_20 = 288'hC2A33FF84C633000C0FFA11898D06335998C667FD08C4C2A33FF84C633000C0FFA1189FF;
defparam spx9_inst_2.INIT_RAM_21 = 288'h06337008CFFA118985C663198C5621D8EC6131880C67630E10198D06335998C667FD08C4;
defparam spx9_inst_2.INIT_RAM_22 = 288'hC63331B8C467FD08C4C2E3318CC007FF08CC66233FF84C663199FF42310000CFFA1189AC;
defparam spx9_inst_2.INIT_RAM_23 = 288'h06335988CFFE13198C667FD08C4C0233FE8462617198C66003FFFFFFA118980C66B3198C;
defparam spx9_inst_2.INIT_RAM_24 = 288'h62003FF84D2B319ACC467FF098CC6333580C668031A0C66B3318CCFFE134ACC6680181AC;
defparam spx9_inst_2.INIT_RAM_25 = 288'h423130B8CC633001FFFFA118980C66B3198CC63331B8C467FD08C4C2E3318CC00033FE84;
defparam spx9_inst_2.INIT_RAM_26 = 288'h3B1D8C2631018CEC61C2030000CFFA1189FF4231001FFFFE0319ACC663318CCC6E3119FF;
defparam spx9_inst_2.INIT_RAM_27 = 288'hC663198C4FFE13198C66313FF84C66319800067FD08C4FF813FE04C68319BFF423118AC4;
defparam spx9_inst_2.INIT_RAM_28 = 288'h3B1D8C2631018CEC61C2033FF8466333598C1633599ACC60B19ACCC6333FF8466313FF84;
defparam spx9_inst_2.INIT_RAM_29 = 288'h319D8C384067FF09ACC66319AC4FFE13198C6600019FF42313FF8D06337FE84623158AC4;
defparam spx9_inst_2.INIT_RAM_2A = 288'hFFB13580C66B13FF84C663198C4FFE13198C6600019FF423131A0C66B1588763B184C620;
defparam spx9_inst_2.INIT_RAM_2B = 288'h3B187080CFFA118800FFA1188C5FFB13580C66803FE8462317FEC4D60319A00FFA1188C5;
defparam spx9_inst_2.INIT_RAM_2C = 288'hFFFFD88C4FFE13198C6600019FF42313FE04C68319BFFFFA1188C562B10EC763098C4063;
defparam spx9_inst_2.INIT_RAM_2D = 288'h3098C40633B187098C6600019FF423131A0C66E3418CD66230EC763098C40633B187080C;
defparam spx9_inst_2.INIT_RAM_2E = 288'h42313FE846260119FFC26959B8CC633198CD6733F198DC763F18CCFFA1188C5621D8EE76;
defparam spx9_inst_2.INIT_RAM_2F = 288'h6663198CCC6330000CFFA1189AC06337008CFFE134ACDC66319800067FD08C4FFA1189FF;
defparam spx9_inst_2.INIT_RAM_30 = 288'h66331D88CFFE13198C666DC188DFFE13198C66331D88CFFE13198C666DC188DFFE1318CC;
defparam spx9_inst_2.INIT_RAM_31 = 288'hC633198EC467FF098CC63336E0C46FFF098C66331D88CFFE13198C666DC188DFFE13198C;
defparam spx9_inst_2.INIT_RAM_32 = 288'h0633598EC467FF098CC63336E0C46FFF098CC633198EC467FF098CC63336E0C46FFF098C;
defparam spx9_inst_2.INIT_RAM_33 = 288'hFFA1189806633018000663418CDC68319B8D063371A0C66EB018CDC03331A0C66E01998D;
defparam spx9_inst_2.INIT_RAM_34 = 288'hFFE134ACDC66319800FF8130ACC6663198CCC6331998C6633318CC6663198CCC6330000C;
defparam spx9_inst_2.INIT_RAM_35 = 288'h66331D88CFFE13198C666DC188DFFE1318CC6663198CCC6330000CFFA1189AC06337008C;
defparam spx9_inst_2.INIT_RAM_36 = 288'hC633198EC467FF098CC63336E0C46FFF098C66331D88CFFE13198C666DC188DFFE13198C;
defparam spx9_inst_2.INIT_RAM_37 = 288'h0633598EC467FF098CC63336E0C46FFF098CC633198EC467FF098CC63336E0C46FFF098C;
defparam spx9_inst_2.INIT_RAM_38 = 288'hFFA1149806633018000663418CDC68319B8D063371A0C66EB018CDC03331A0C66E01998D;
defparam spx9_inst_2.INIT_RAM_39 = 288'hC263318CCC0233FF84D2B37198C6600018CCC6331998C6633318CC6663198CCC6330000C;
defparam spx9_inst_2.INIT_RAM_3A = 288'hD60319A000633318CC666319800067FD08A4C0633598CC6733198C67637598C7633589FF;
defparam spx9_inst_2.INIT_RAM_3B = 288'h067FD08A462B198FFF422918AC663B3198CC6633198CC6633198CC667FC0985667FD08A4;
defparam spx9_inst_2.INIT_RAM_3C = 288'h62313FF84C66319800067FD08A4FFE3418CDFFA1148C562B10EC763098C40633B9D8C384;
defparam spx9_inst_2.INIT_RAM_3D = 288'h62B10EC763098C40633B1870800FF8130ACCFFE1198C5621D8EC6131880C67630E1019FF;
defparam spx9_inst_2.INIT_RAM_3E = 288'h66233FF84C663198CC467FF098CC6331988CFFE13198C667FD08A400033FE84526B018CD;
defparam spx9_inst_2.INIT_RAM_3F = 288'h3B184C620319D8C384067FF09A566337FE845261599FF422930ACC66633598C6663718CC;

SPX9 spx9_inst_3 (
    .DO({spx9_inst_3_dout_w[26:0],spx9_inst_3_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_3.READ_MODE = 1'b0;
defparam spx9_inst_3.WRITE_MODE = 2'b01;
defparam spx9_inst_3.BIT_WIDTH = 9;
defparam spx9_inst_3.BLK_SEL = 3'b011;
defparam spx9_inst_3.RESET_MODE = "SYNC";
defparam spx9_inst_3.INIT_RAM_00 = 288'h66637598C76637198C66313FF84C663198C4FFE13198C6600019FF42293580C66B158876;
defparam spx9_inst_3.INIT_RAM_01 = 288'hFFE13198C6631588763B184C620319D8C384067FD08A4C2B31988CFFE1198CCD6633198C;
defparam spx9_inst_3.INIT_RAM_02 = 288'hC0331988CFFE13198C6633018000663418CDC68319B8D063371A0C66B13FF84C663198C4;
defparam spx9_inst_3.INIT_RAM_03 = 288'hC60331BADC60331B8C066379ACDC60331CCC006361B8C0600019FF42293FE84527FD08A4;
defparam spx9_inst_3.INIT_RAM_04 = 288'h3098C40633B187080CC6F375AEDC60331D8C0667D98CCC6333FE845261719AC06335998C;
defparam spx9_inst_3.INIT_RAM_05 = 288'hD60319B8D063371BCD068331C0CC033189FFC263318CC00033FE84526B018CD62B10EC76;
defparam spx9_inst_3.INIT_RAM_06 = 288'hF68331C0C006379A0D06638198DE6EB7DA0CC7030018DE6EB7DA0CC703001AC0633700CC;
defparam spx9_inst_3.INIT_RAM_07 = 288'hC6030EC763098C40633B187080CC6837180C00033FE8452000018DE6834198E066379BAD;
defparam spx9_inst_3.INIT_RAM_08 = 288'h6680198CCC683419FF42293FF8DE683419AEC67B19A00660331A0DC60331A0DC60331A0D;
defparam spx9_inst_3.INIT_RAM_09 = 288'h6633000CC066B018CD66631998DE683419AEC67B19B8D66E3198CCC63331BAD66637580C;
defparam spx9_inst_3.INIT_RAM_0A = 288'h3098C40633B187080CD60319ACCC63331ACDC6331998C667FD08A4D6633980C676359800;
defparam spx9_inst_3.INIT_RAM_0B = 288'h4229001FFC26B018CD007FE09AC0633589FFC263318CC00033FE84526B018CD62B10EC76;
defparam spx9_inst_3.INIT_RAM_0C = 288'h30E1001FF422930ACC66233FF8D068331A0D0631588763B184C620319D8C3840600019FF;
defparam spx9_inst_3.INIT_RAM_0D = 288'h6600180CC067FD08A460313FF84C66319800067FD08A4D60319AC5621D8EC6131880C676;
defparam spx9_inst_3.INIT_RAM_0E = 288'hFFE118A06D63319BFF422931A0C66B3318CCC6EB79BAC663371DAC066B598CD00301998C;
defparam spx9_inst_3.INIT_RAM_0F = 288'hC66319800067FD08A4D60319AC5621D8EC6131880C67630E1019FF4229358CC66B3318CC;
defparam spx9_inst_3.INIT_RAM_10 = 288'hE60339CCC6763758CC6680181FFC23140DAC66335998C6600180CC067FD08A460313FF84;
defparam spx9_inst_3.INIT_RAM_11 = 288'h66B3318CCFFA11498D06335998C66003FE84527170DAC066B598CDC763358CC66EB3198C;
defparam spx9_inst_3.INIT_RAM_12 = 288'h52313FF84C66319800067FD08A4D60319AC5621D8EC6131880C67630E1019FF4229358CC;
defparam spx9_inst_3.INIT_RAM_13 = 288'h66233FF8D068331A0D0630180C5621D8EC6131880C67630E1019FFC26B018CDFFB13FE84;
defparam spx9_inst_3.INIT_RAM_14 = 288'h663371DAC066B598CD00301998C6600180CC067FD08A4FFE13580C66FFD89FF422930ACC;
defparam spx9_inst_3.INIT_RAM_15 = 288'hFFA1149FF4229358CC66B3318CCFFA1149FFC23140DAC663371A0C66B3318CCC6EB79BAC;
defparam spx9_inst_3.INIT_RAM_16 = 288'hC66B198CDD663319CC0673998CEC6EB198CD00303FF846281B58CC66B3318CC00301980C;
defparam spx9_inst_3.INIT_RAM_17 = 288'hC2033FE84526B198CD6663199FF422931A0C66B3318CC007FD08A4E2E1B580CD6B319B8E;
defparam spx9_inst_3.INIT_RAM_18 = 288'hC2B31980C66031980C6663019FFC2333FF84060140DFFC20300A063B1D8C2631018CEC61;
defparam spx9_inst_3.INIT_RAM_19 = 288'h319DB080C6031588763B18C40633B187080CFFB1588763B184C620319D8C384007FF080C;
defparam spx9_inst_3.INIT_RAM_1A = 288'hC6EB018CDC76B018CD00303584C66B3318CCC06B018CD00303FE845231588763B184C620;
defparam spx9_inst_3.INIT_RAM_1B = 288'h422918BC6C3E33580C66E3B580C66EB319CC0633B1BAC0633400C0D61319ACCC633359CC;
defparam spx9_inst_3.INIT_RAM_1C = 288'h3B18401FFC20300BFF422900AC6531D8EC6131880C67630E101980066B098CD6663199FF;
defparam spx9_inst_3.INIT_RAM_1D = 288'h02FFD08A402B194C763B184C620319D8C200FFE101805FFA11480563298EC763098C4063;
defparam spx9_inst_3.INIT_RAM_1E = 288'h531D8EC6131880C67630803FF8406017FE84420158CA63B1D8C2631018CEC61007FF080C;
defparam spx9_inst_3.INIT_RAM_1F = 288'h319D8C200FFE101805FFA11080563298EC763098C40633B18401FFC20300BFF422100AC6;
defparam spx9_inst_3.INIT_RAM_20 = 288'h06017FE84420158CA63B1D8C2631018CEC61007FF080C02FFD088402B194C763B184C620;
defparam spx9_inst_3.INIT_RAM_21 = 288'h63298EC763098C40633B18401FFC20300BFF422100AC6531D8EC6131880C67630803FF84;
defparam spx9_inst_3.INIT_RAM_22 = 288'h1018CEC61007FF080C02FFD088402B194C763B184C620319D8C200FFE101805FFA110805;
defparam spx9_inst_3.INIT_RAM_23 = 288'hC20304BFF422100AC6531D8EC6131880C67630803FF8406017FE84420158CA63B1D8C263;
defparam spx9_inst_3.INIT_RAM_24 = 288'h02B190C763B184C620319D8C200FFE101845FFA11080563298EC763098C40633B18401FF;
defparam spx9_inst_3.INIT_RAM_25 = 288'h31880C67630803FF8406417FE84420158C863B1D8C2631018CEC61007FF080C42FFD0884;
defparam spx9_inst_3.INIT_RAM_26 = 288'hFFE101805FFA11080563218EC763098C40633B18401FFC20300BFF422100AC6431D8EC61;
defparam spx9_inst_3.INIT_RAM_27 = 288'h420158C863B1D8C2631018CEC61007FF080C02FFD088402B190C763B184C620319D8C200;
defparam spx9_inst_3.INIT_RAM_28 = 288'h3098C40633B18401FFC20300BFF422100AC6431D8EC6131880C67630803FF8406017FE84;
defparam spx9_inst_3.INIT_RAM_29 = 288'h007FF080C02FFD088402B190C763B184C620319D8C200FFE101805FFA11080563218EC76;
defparam spx9_inst_3.INIT_RAM_2A = 288'h422100AC6431D8EC6131880C67630803FF8406017FE84420158C863B1D8C2631018CEC61;
defparam spx9_inst_3.INIT_RAM_2B = 288'h3B184C620319D8C200FFE101805FFA11080563218EC763098C40633B18401FFC20300BFF;
defparam spx9_inst_3.INIT_RAM_2C = 288'h30803FF8406017FE84420158C863B1D8C2631018CEC61007FF080C02FFD088402B190C76;
defparam spx9_inst_3.INIT_RAM_2D = 288'hFFA11080563218EC763098C40633B18401FFC20300BFF422100AC6431D8EC6131880C676;
defparam spx9_inst_3.INIT_RAM_2E = 288'h3B1D8C2631018CEC61007FF080C02FFD088402B190C763B184C620319D8C200FFE101805;
defparam spx9_inst_3.INIT_RAM_2F = 288'hC663019FF422100AC6436341B8C061D8EC6131880C67630803FF8406017FE84420158C86;
defparam spx9_inst_3.INIT_RAM_30 = 288'h308031A0C66B3318CCC0E33598C666B51B80C66B198CD0030000CCD63319ACCC663018CC;
defparam spx9_inst_3.INIT_RAM_31 = 288'h66633198CC663118763B184C620319D8C200FFB33198C066341B8C061D8EC6131880C676;
defparam spx9_inst_3.INIT_RAM_32 = 288'hC66341B8C061D8EC631018CEC61007FD0884C2B331A0DC62331A0DC6031998CC6633188C;
defparam spx9_inst_3.INIT_RAM_33 = 288'hC62331ACCC68319B8DE6837180CC763018CCC6633198C061D8EC6131880C67600333198C;
defparam spx9_inst_3.INIT_RAM_34 = 288'h3B184C620319D8C200000031BCDD6BB7180CC763019FF422100180C6033FE844260319AC;
defparam spx9_inst_3.INIT_RAM_35 = 288'hC6837180CFFA11098566333190CC063199FF42213FE04C0233FE04C063198CCC66301876;
defparam spx9_inst_3.INIT_RAM_36 = 288'hFF9D8EC6131880C676308031A0DC60331A0DC6033FF84667FD0884C2B31998C0660318CC;
defparam spx9_inst_3.INIT_RAM_37 = 288'h0049609AC5DA6818ED002E530F79B984F67A3C9E0EE63000000020319D8C200FFFFD0884;
defparam spx9_inst_3.INIT_RAM_38 = 288'h32180C0E03C9E0F278301B3188C363DC1820319ECF4793C1DECB4430A0001258201C0C80;
defparam spx9_inst_3.INIT_RAM_39 = 288'h003B0186532001CAC40381BFE8C3D9E8D8001018CF67A3C9E0EF65A2184F67AC01B10000;
defparam spx9_inst_3.INIT_RAM_3A = 288'h082139B8CD6F839BACE623F1A0D4263100A402A39580D4C2DF60613C1DC1A63007FD180C;
defparam spx9_inst_3.INIT_RAM_3B = 288'h1074C61CCF8903DFADC614B638E000001E120A07FDFADC6297182EC884365D10003C1C05;
defparam spx9_inst_3.INIT_RAM_3C = 288'h31E94F077821875B184694A31B70B9615AAC0C24B018C2FFBF5B8C37250A5B1D6E335D8C;
defparam spx9_inst_3.INIT_RAM_3D = 288'h3984FFFACC21379DB039F48261FF8EC35A2F000481FE00787F9C0DC6741401F568416020;
defparam spx9_inst_3.INIT_RAM_3E = 288'h430014E861018F4A783BC115A9830801CF060029D0DFF29249180CFF8332620186C7FFD3;
defparam spx9_inst_3.INIT_RAM_3F = 288'h426B55A0CD76B41BAE0603B5A0D56033008C00003FE0F09F4BFEA5FF8315BFF56A6000A7;

SPX9 spx9_inst_4 (
    .DO({spx9_inst_4_dout_w[26:0],spx9_inst_4_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[17:9]})
);

defparam spx9_inst_4.READ_MODE = 1'b0;
defparam spx9_inst_4.WRITE_MODE = 2'b01;
defparam spx9_inst_4.BIT_WIDTH = 9;
defparam spx9_inst_4.BLK_SEL = 3'b000;
defparam spx9_inst_4.RESET_MODE = "SYNC";
defparam spx9_inst_4.INIT_RAM_00 = 288'hFF7C411FE000210018007F01000040000000007A0349000000000800868021A940002080;
defparam spx9_inst_4.INIT_RAM_01 = 288'h0000000000000000000000000000000000000000000000010000EE7C000001090080A122;
defparam spx9_inst_4.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam spx9_inst_4.INIT_RAM_20 = 288'h0B1002C200B0402C08195E0152194CC67341A4D46B361B4EE783C9E8F67C3E9F8FE40062;
defparam spx9_inst_4.INIT_RAM_21 = 288'hB0DA773C1E4F47B3E1F4FC7F200013580C80055681D86091E82C600D0783DFE0B0002D00;
defparam spx9_inst_4.INIT_RAM_22 = 288'hEB804000CEF1682C001C040017000003F000007A3F440057A0386290CA66339A0D26A359;
defparam spx9_inst_4.INIT_RAM_23 = 288'hECF87D3F1FC800C400FD20015E8F780801E8FD10015E8090010000040039614F6FFBF048;
defparam spx9_inst_4.INIT_RAM_24 = 288'h011E3D7008418803118CC8653319CD069351ACD86D371BCE071391CCE8753B1DCF0793D1;
defparam spx9_inst_4.INIT_RAM_25 = 288'h9CD069351ACD86D371BCE071391CCE8753B1DCF0793D1ECF87D3F1FC803130800100F1FC;
defparam spx9_inst_4.INIT_RAM_26 = 288'hEB8980418EBED46DD7EC80373C1ECF276BA9406E4C058D0000C4000418A13118CC865331;
defparam spx9_inst_4.INIT_RAM_27 = 288'h2C68000602C00001D9DCF203DD7EB80BAFD94C76731C9D4F64B1D90C7078398E481B9242;
defparam spx9_inst_4.INIT_RAM_28 = 288'h007000818ECEE7CE16ECFE011C00179C01EAECEC7B202EC81001E70C7677214ECEC77260;
defparam spx9_inst_4.INIT_RAM_29 = 288'hECEC772602C68000602C00001C00206373FED8F9FF002E000BCE00F276501FED8F6405D9;
defparam spx9_inst_4.INIT_RAM_2A = 288'hF3863B3B9007000818E8EE7CFF80170005E7000D3A3EA03767B202EC81001E70C7677214;
defparam spx9_inst_4.INIT_RAM_2B = 288'h00773A3B1E880BA200E001031D1DCF9FF002E000BCE001172BB3B1E880BA3D9017640800;
defparam spx9_inst_4.INIT_RAM_2C = 288'hF3F0015E710063C00010060000AE016BBDE7E002BCE0AE000BCFC00579C4018F0000C058;
defparam spx9_inst_4.INIT_RAM_2D = 288'h200C07080EDEFD1680027673BD90576480301C70000200C00015C01079F800AF382B8002;
defparam spx9_inst_4.INIT_RAM_2E = 288'h180E0017B23A0005D9ACF5FB20CEC9006038E000040100C003F40240744002008063C000;
defparam spx9_inst_4.INIT_RAM_2F = 288'h30140B1A000100603840003B34B0BA0009D90FA0011D998F7FBBDBECC8080301C7000040;
defparam spx9_inst_4.INIT_RAM_30 = 288'h00180A0580053E03CD40023B2DFBCF6F81B9DC94373DDE06E77250DCF7F81B9ECEC3B3B9;
defparam spx9_inst_4.INIT_RAM_31 = 288'hD4E050008ECA4E5BDBE06E77250DCF7781B9DC94373DFE06E7B204ECEA763B930140B1A0;
defparam spx9_inst_4.INIT_RAM_32 = 288'hDCEE4A1B9EEF0373B9286E7BFC0DCF640DD9D4EC7726028163400030140B0007EABFE7B1;
defparam spx9_inst_4.INIT_RAM_33 = 288'h9000080301C0023DE84077FBE80200C071C000180A0580017F47B1D4CC50008EC90FB7C0;
defparam spx9_inst_4.INIT_RAM_34 = 288'h94D8035E1EC8BA00046C7265228ECF267206E196B92989C83A721290C8653319CB81A0D8;
defparam spx9_inst_4.INIT_RAM_35 = 288'h0970782800258031E1FF7441DD9E88EBA298CD76A31D9ECCC7B1C9EC80BB3C98001135C9;
defparam spx9_inst_4.INIT_RAM_36 = 288'h03053BE18DC980A058D0001C0D06C20101C6E8F47FDD1A5A0380AEE070415C030703820C;
defparam spx9_inst_4.INIT_RAM_37 = 288'h208E46229108642209CCA00E078A0000C0502C20101E2EFF7C01B9DC80B73194077E3E1A;
defparam spx9_inst_4.INIT_RAM_38 = 288'h0074400000C3C00044AB29B6C000C66405D9E480AE44AE3F1C0018CCF6731D9E8EE773C8;
defparam spx9_inst_4.INIT_RAM_39 = 288'hECF4411D144A03921440003A334EC80BB3D1047450E80E0003A34CEC80BB3D104746DA80;
defparam spx9_inst_4.INIT_RAM_3A = 288'hE8B83B202ECF4411D128A03921040003A2FCEC80BB3D104744DA80E48500400E8C63B202;
defparam spx9_inst_4.INIT_RAM_3B = 288'hEC80BB3E9252A3B202ECF4411D10CA03922040003A2C4EC80BB3D1047446A80E48110000;
defparam spx9_inst_4.INIT_RAM_3C = 288'h000633202ECBB0C0000C66405D9EC80BB3C90C6800018CC80BB2180A7243DC9EC80BB29C;
defparam spx9_inst_4.INIT_RAM_3D = 288'h390003199017655C60000633202ECF6405D9E486340000C66405D90C053921EE4B779472;
defparam spx9_inst_4.INIT_RAM_3E = 288'hDC980B1A000300E07840200C4000C667B3D9017668E80E3D3434060A71C2400AD9293FCA;
defparam spx9_inst_4.INIT_RAM_3F = 288'h066E405B9036E780FEE001B7202DC80015B9026537206DCF013100E001B7206036E7A3DF;

SPX9 spx9_inst_5 (
    .DO({spx9_inst_5_dout_w[26:0],spx9_inst_5_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[17:9]})
);

defparam spx9_inst_5.READ_MODE = 1'b0;
defparam spx9_inst_5.WRITE_MODE = 2'b01;
defparam spx9_inst_5.BIT_WIDTH = 9;
defparam spx9_inst_5.BLK_SEL = 3'b001;
defparam spx9_inst_5.RESET_MODE = "SYNC";
defparam spx9_inst_5.INIT_RAM_00 = 288'h000204018F0000803800003AFD9FC103800AEC803AE80EC90071C000180B000EF8037204;
defparam spx9_inst_5.INIT_RAM_01 = 288'h1C70000200C001100210063C00010060008210063C0001006000000408031E0000803000;
defparam spx9_inst_5.INIT_RAM_02 = 288'hE8863D7D10C764B1FE0780021EBE8F64A1B91A6E772602C68000401C001040641767B240;
defparam spx9_inst_5.INIT_RAM_03 = 288'h0077C5C00047A37E803016340003016000002D3F811EB00023D6120040011EB00023D600;
defparam spx9_inst_5.INIT_RAM_04 = 288'hEF80373B9016E77280EFEFC34060A77C31B930140B1A000180B000006FFD1F8020105DDF;
defparam spx9_inst_5.INIT_RAM_05 = 288'hE4CA451D9E4CE40D7B2D7253139074E4252190CA6633970341B12000180A05840203C5DF;
defparam spx9_inst_5.INIT_RAM_06 = 288'hE883BB3D11D745319AED463B3D998F6393D90176793000226B9329B006BC3D91740008D8;
defparam spx9_inst_5.INIT_RAM_07 = 288'h00381A0D8402038DD1E8FFBA303407015DC0E082B8060E07041812E0F050004B0063C3FE;
defparam spx9_inst_5.INIT_RAM_08 = 288'hCC80BB3C9015C895BFDF8003199ECF03B3D1D8EC790411C8C452210C8441399401C0F140;
defparam spx9_inst_5.INIT_RAM_09 = 288'h01767A208E89DD01C00074699D901767A208E8AF50000E88000018940008956536D80018;
defparam spx9_inst_5.INIT_RAM_0A = 288'h00745F9D901767A208E8A9501C90A00801D18C76405D9E8823A2C14072428800074669D9;
defparam spx9_inst_5.INIT_RAM_0B = 288'h4072440800074589D901767A208E89B501C90220001D17076405D9E8823A289407242080;
defparam spx9_inst_5.INIT_RAM_0C = 288'h017679218D00003199017643014E487B93D90176539D901767B24A5476405D9E8823A251;
defparam spx9_inst_5.INIT_RAM_0D = 288'hEC80BB3C90C6800018CC80BB2180A7243DC96EF28E4000C66405D9761800018CC80BB3D9;
defparam spx9_inst_5.INIT_RAM_0E = 288'h2D07BB226ECCDD01BF9E8680C14DF848014B2527F9472000633202ECAB8C0000C66405D9;
defparam spx9_inst_5.INIT_RAM_0F = 288'h200E38000601C0F080400E80018CCF67B202ECFCB83FEE080000000002B82660006A0004;
defparam spx9_inst_5.INIT_RAM_10 = 288'hECF6480301C70000200C002BC2010063C00010060015E1008031E0001007080ECF6461D9;
defparam spx9_inst_5.INIT_RAM_11 = 288'h0A26001B9046E41C00DC8237208DCA0333B930140B1A000100603800003B280DA823B200;
defparam spx9_inst_5.INIT_RAM_12 = 288'hECF673E80E482B0680E4D97A3C9ECEE4C0502C6800060281610018046E531D9006E7B3FE;
defparam spx9_inst_5.INIT_RAM_13 = 288'h400610000ECF6480301C7000040180E001BD4011BB3D9200C071C000180A0580057FE9B9;
defparam spx9_inst_5.INIT_RAM_14 = 288'h03003B202EC843A3D9200E38000200C07000E7A0031D0ECF6480301C7000040180E0019D;
defparam spx9_inst_5.INIT_RAM_15 = 288'hEC80031EBE8F6772602C68000401C2013000E8F47FDD140003B3E60074405D1007644480;
defparam spx9_inst_5.INIT_RAM_16 = 288'hE881373C01F700C1D1036E7803EE076411B9E007B804AEC82B73C07F700A5D9E880021EB;
defparam spx9_inst_5.INIT_RAM_17 = 288'hEC82005D904023B2080C023B3D9200E38000301600000DCF00FDC02474405B9E01FB8054;
defparam spx9_inst_5.INIT_RAM_18 = 288'h3C003B2982A70200046C1E005D93070200046C0C009D900003D606017641006EC8207C06;
defparam spx9_inst_5.INIT_RAM_19 = 288'h1F01BB2982570200046C06811D92902BB200087AD35C080011B4C8067653048E040008D8;
defparam spx9_inst_5.INIT_RAM_1A = 288'hD000080301C00263D103307A208EFF7FA280200C071C00010070000000011EB00063D698;
defparam spx9_inst_5.INIT_RAM_1B = 288'h1A20139EB40663B202407AC90802E7AD0018CC7640480F586363D9DC8D07DB9D8EE4C058;
defparam spx9_inst_5.INIT_RAM_1C = 288'h3016340003016000A04E7AD0198EC80941EB0A280B9EB4006331D901283D618D8F6781B9;
defparam spx9_inst_5.INIT_RAM_1D = 288'hE06E468884E7AD0198EC80911EB24220B9EB4006331D901223D618D8F6772341F6E763B9;
defparam spx9_inst_5.INIT_RAM_1E = 288'h007A84018F0000C058002A139EB40663B202547AC28A82E7AD0018CC76404A8F586363D9;
defparam spx9_inst_5.INIT_RAM_1F = 288'h047AC0008F5800B5FEFF823D600047AD4018D8F6763B9301634000100600000E0023D5C0;
defparam spx9_inst_5.INIT_RAM_20 = 288'hD88237200DCA6001B1006E421B94C0036210DC84021B92C06001B1086E42808D88013400;
defparam spx9_inst_5.INIT_RAM_21 = 288'h0C6E53000D88637208DC9603000D88237212046E53000D88237212010436208DC9603000;
defparam spx9_inst_5.INIT_RAM_22 = 288'hE0000803800063B210017641002EC803B3D9200E38000301600000DC9603000D88037212;
defparam spx9_inst_5.INIT_RAM_23 = 288'h200E000604D767D6600C764D154AD7AFB2401C70000401C00031D94C74431D9E8F648038;
defparam spx9_inst_5.INIT_RAM_24 = 288'hECC00089AE88036204206E7A2003D76763B930140B1A000080300034552B5EB10063C000;
defparam spx9_inst_5.INIT_RAM_25 = 288'hDC82019B1026E7809880701300ED8F01300CD88236202DCF00A1D9006E781D9ECFF889D9;
defparam spx9_inst_5.INIT_RAM_26 = 288'h077641804EC828A9D904103B200A0007B3D9200E3800030140B0008F7A41DB9056C41008;
defparam spx9_inst_5.INIT_RAM_27 = 288'hE0000803800023B3C02C5FB8008EC84811D9E02038008EC84BA3D1EC90071C0001007000;
defparam spx9_inst_5.INIT_RAM_28 = 288'hE072781D14D76793D1EC9006038E000080301C0001020F481BAFD961767AE80EC9006038;
defparam spx9_inst_5.INIT_RAM_29 = 288'h8400101D7EB80BAE14EA993B3D54075D0080EC9006038E000080301C00011D9E01038098;
defparam spx9_inst_5.INIT_RAM_2A = 288'h046E411DF046E772602C6800040180E00008907A40DD7ECD4DE0004075FAE58FE75C2967;
defparam spx9_inst_5.INIT_RAM_2B = 288'h281634000301600008DCF0011C0046E42008EFF7C11B9DC980B1A000180B000FB013BFDF;
defparam spx9_inst_5.INIT_RAM_2C = 288'hE0023D375F4C8FD2804077D7AC80020101BBEFF7E81C0E013B7BBDFF6F77680DEA010060;
defparam spx9_inst_5.INIT_RAM_2D = 288'h40FA501BB38FA000081770011E9A3FA53BE9407037A8F4400101BDDEFFB7A9F50000102E;
defparam spx9_inst_5.INIT_RAM_2E = 288'hE013B7BBDFF6F77A8030140B1A000180A05800447D231F4808AB78000205DC0047A657E9;
defparam spx9_inst_5.INIT_RAM_2F = 288'hDEEF7FDBDF89E00080DEFED1000040BB8008F4B47D27FF4A0101DF0CB200080EFF7E81C0;
defparam spx9_inst_5.INIT_RAM_30 = 288'hF484101AFAC000102EE0023D285F48CFD2800177F9BD0000205DC0047A547E9FCFA501C0;
defparam spx9_inst_5.INIT_RAM_31 = 288'h007D005D9EC80021EC057640010F60000010F610071C000180A05840777BA06F49A7D3E7;
defparam spx9_inst_5.INIT_RAM_32 = 288'hD48036208F6000B5FEFFEE7D9F401767B200087B015D900043D9A9D8EE4C058D00008038;
defparam spx9_inst_5.INIT_RAM_33 = 288'h2C7F8005E02765306001764E000ECF648038E0000C058000000410F60280006087B01802;
defparam spx9_inst_5.INIT_RAM_34 = 288'h4C161806C01764E000ECF648038E000080380000021EB4C07811D94C16000002801BB298;
defparam spx9_inst_5.INIT_RAM_35 = 288'h0017809D930003B3D9200E38000200E000000C7AD3408ECA6000500376530581F98009D9;
defparam spx9_inst_5.INIT_RAM_36 = 288'h01043B298021081DD94C7F8900CECA6000500576530002B023B2982C000B006ECA60B1FE;
defparam spx9_inst_5.INIT_RAM_37 = 288'h200E000002D7F811EB00023D6120000011EB00023D612ECF648038E0000803800003D698;
defparam spx9_inst_5.INIT_RAM_38 = 288'h0006201EB40113BBDD4010071C0001007080E07FB80000C203D68022777BA80200E38000;
defparam spx9_inst_5.INIT_RAM_39 = 288'hE000040180000005EB007AC4018F000040180000009EB007AC4018F0000803840703FDC0;
defparam spx9_inst_5.INIT_RAM_3A = 288'h1C70000401C000009C0D203D6802277D0070EEFF80018407AD0044EFF7501DF402008038;
defparam spx9_inst_5.INIT_RAM_3B = 288'h281634000200E000004C06901EB40113BFFE0006201EB40113BE8038777BA80EFA010040;
defparam spx9_inst_5.INIT_RAM_3C = 288'hE9883A2A0CFA0100703C60000602816001EA0B777BA02EEEA50080DFF03BA14EEEFD0060;
defparam spx9_inst_5.INIT_RAM_3D = 288'hDA81B6606D8EBC0DAD016A7FDBF4070793FEE38438A10E1F040D8F40747B202EB80BAA02;
defparam spx9_inst_5.INIT_RAM_3E = 288'h401B501C0EC87BB2A048262C000401C0F0001880AC280CFFE80400F5801BBE3406A773B7;
defparam spx9_inst_5.INIT_RAM_3F = 288'hF205BB3D901767EB68002032018F0913B21AEC82C1000F005BB3D9017672018F0913B280;

SPX9 spx9_inst_6 (
    .DO({spx9_inst_6_dout_w[26:0],spx9_inst_6_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[17:9]})
);

defparam spx9_inst_6.READ_MODE = 1'b0;
defparam spx9_inst_6.WRITE_MODE = 2'b01;
defparam spx9_inst_6.BIT_WIDTH = 9;
defparam spx9_inst_6.BLK_SEL = 3'b010;
defparam spx9_inst_6.RESET_MODE = "SYNC";
defparam spx9_inst_6.INIT_RAM_00 = 288'h0C7B40008EC843DA00047B401EDEC90071C00028120980074E70004075FAE1EE000011EB;
defparam spx9_inst_6.INIT_RAM_01 = 288'hF68C3B200F680135ED1076401ED0070005EAE0003D41014764009AF68A3B200F680021D9;
defparam spx9_inst_6.INIT_RAM_02 = 288'hEC8420001EC820FC00EC88011D914013B2300176400003D767B2401C70000401C000009A;
defparam spx9_inst_6.INIT_RAM_03 = 288'h0E767B2401C70000401C00001FCF6803DA0C0000BDA00F683BB3D9200E38000200E00018;
defparam spx9_inst_6.INIT_RAM_04 = 288'h2C68000401C00001C02D7F3D5C0007A801FAF6803DA1C0070005EAE0003D400027B401ED;
defparam spx9_inst_6.INIT_RAM_05 = 288'hF57000006F500135D9F6803DBD9200E380003016101D9EC813B202041637200F6F677260;
defparam spx9_inst_6.INIT_RAM_06 = 288'hEC90071C000100603800032D1FF4077C0002C87FFBE80200C071C0001007000007000406;
defparam spx9_inst_6.INIT_RAM_07 = 288'hEC88811D91076441D901083B218EC81811D90C76431D901063B200EB86831D900767AE80;
defparam spx9_inst_6.INIT_RAM_08 = 288'h281634000200E10000E8F648038E0000803800043B2060476421D9087640410EC883B208;
defparam spx9_inst_6.INIT_RAM_09 = 288'h0076405D9B88E00080400003048ECA600002EC88BB38F48001AC48026E41402DCEC77260;
defparam spx9_inst_6.INIT_RAM_0A = 288'h2476680001A200F3D1400003048ECE600050ECF4411B14E729009BE800100000C123B228;
defparam spx9_inst_6.INIT_RAM_0B = 288'h00200001824764C000EC80BB22080A40008040200301824765C0000806091D9880000018;
defparam spx9_inst_6.INIT_RAM_0C = 288'hC0000C0502C2010000022EFA0000530F60000920023A8002000018247640000CE2005208;
defparam spx9_inst_6.INIT_RAM_0D = 288'hE880000000002BA266002561000F9767FDD9000000000057671C1C0002811E881A00E078;
defparam spx9_inst_6.INIT_RAM_0E = 288'h29201002040200000830003E5C9FF72400000000015C933000DE88006874298007CBA3FE;
defparam spx9_inst_6.INIT_RAM_0F = 288'h056E4CC0005CA00080C4E2421F2E0FFB820000000000AE09980031D400333914110F3280;
defparam spx9_inst_6.INIT_RAM_10 = 288'hE403A0202017CB63FED880000000002B63C80766D4A28012AC0402F96E7FDB9000000000;
defparam spx9_inst_6.INIT_RAM_11 = 288'hDC82005B9D8EE4C0502C68000200C20100200C7838AE301203E5A9FF6A400000000015A9;
defparam spx9_inst_6.INIT_RAM_12 = 288'hEC8401DD917767A280B32000010D8843A2020401373C9BF2000008D8980055F880001806;
defparam spx9_inst_6.INIT_RAM_13 = 288'hDC980A058D0000C0502C20101D0E8F67B202ECC2C3000407000018E4F663A480020031C9;
defparam spx9_inst_6.INIT_RAM_14 = 288'hECF4500DC4000021B1087440408026E792F44000011B133009AB50000300DB90400B73B1;
defparam spx9_inst_6.INIT_RAM_15 = 288'h2C20101CAE8F67B202EC9EC70004000031C940113B28F380010018E4A0089D90A01BB234;
defparam spx9_inst_6.INIT_RAM_16 = 288'hEBF67AE802F2000010D8F64D4800002362240112F10000601B73B1DC980A058D0000C050;
defparam spx9_inst_6.INIT_RAM_17 = 288'h0B2000010D8F6444800002362220100D50000601B73B1DC980A058D0000C0502C2010000;
defparam spx9_inst_6.INIT_RAM_18 = 288'hE481018B00000B720C7800005B91018001B9ECEE4C0502C680006028161008000747B3D1;
defparam spx9_inst_6.INIT_RAM_19 = 288'hE0A18C410E882841D137053A3C10006393B95574429C95974421C901030C000DC86BA220;
defparam spx9_inst_6.INIT_RAM_1A = 288'h467043080E089BB3520C70431D1EC84999C10C3038242ECE8031C10C747B21239704305E;
defparam spx9_inst_6.INIT_RAM_1B = 288'h74AC00008ECE8031C10C747B212E0983A21A2F704502A88C80000AECE4831C10C747B212;
defparam spx9_inst_6.INIT_RAM_1C = 288'h000236232012CC00000601B73B1DC980A058D0000C0502C203B3500006393B9E480B9200;
defparam spx9_inst_6.INIT_RAM_1D = 288'hB800080301C700006028161008040EA00127ECF44048FD40020FD163A000010D8F65A680;
defparam spx9_inst_6.INIT_RAM_1E = 288'h0C203D6802276461D91CD20003F9C00100000C7AC9B48002000010F596EB00040003D667;
defparam spx9_inst_6.INIT_RAM_1F = 288'h3800080301C7000040180E10080E705BB3D9017641AD80076500800006201EB40113B200;
defparam spx9_inst_6.INIT_RAM_20 = 288'h40203DE80E076435D9DC9A001E40B767B202ECF2D400040203E280E076435D9F0BA001E7;
defparam spx9_inst_6.INIT_RAM_21 = 288'h036E45C805AD6000800002363B1DC980A058D000080301C20101E40B767B202ECE8C0000;
defparam spx9_inst_6.INIT_RAM_22 = 288'h026E78002401DD80004000011B18322501DDEEA02F680000436357980024802B0CA0000C;
defparam spx9_inst_6.INIT_RAM_23 = 288'h036E7B6808FA000010D8BEC4000312009238002000008D8B61B3978C9A0000EE01638002;
defparam spx9_inst_6.INIT_RAM_24 = 288'h001C28A804077FB7DF403A500000C6C43808DCA43D816EFF7C05DFB8A0101DFED84BBE1E;
defparam spx9_inst_6.INIT_RAM_25 = 288'h340010000046C474DF3CA40000CE01638002026E780024075DD0004000011B1340094AE8;
defparam spx9_inst_6.INIT_RAM_26 = 288'h50241316000180A058402000802208000047FC000245DEF8238058E000809B9E000901AB;
defparam spx9_inst_6.INIT_RAM_27 = 288'h00062E3D10FA000010B8F64568000022E24E0102CF0008FA01F2800A01AF21F48002E379;
defparam spx9_inst_6.INIT_RAM_28 = 288'h30140B1A000281209840203EE80C8E8430003D72732183F003A3B1227650680C8F242680;
defparam spx9_inst_6.INIT_RAM_29 = 288'h30140B080400250018F828BB3D9D7A000008D8870058F90000120E016E73B18006E763B9;
defparam spx9_inst_6.INIT_RAM_2A = 288'h09F442002ECF46C6800004363D9B7A000008D8978054F280001804DCEC77260281634000;
defparam spx9_inst_6.INIT_RAM_2B = 288'h28161008078B6000087CDC001D113F442006EC8721BB00074437D108013B23090FC001D1;
defparam spx9_inst_6.INIT_RAM_2C = 288'hDAD67B3D96FA000008D885804BF70002E6800800B731F68B8001B9D8EE4C0502C6800060;
defparam spx9_inst_6.INIT_RAM_2D = 288'hAC2800040180E1001EEF81BFC7F080001872EF820BDDFEFA0080301C7000060281610080;
defparam spx9_inst_6.INIT_RAM_2E = 288'h940005B0800079017B40201E200042C613017CBC430100400020002CEC000B15CD829150;
defparam spx9_inst_6.INIT_RAM_2F = 288'hE886163D9082C61C02FCE40000C042E6A080A6A0100F90002163304006F400010DA00027;
defparam spx9_inst_6.INIT_RAM_30 = 288'hECF0432808BA000008EC860288093A000006ECF2432809BA000002EC8602880A3A0001D9;
defparam spx9_inst_6.INIT_RAM_31 = 288'h037476219403650000017443014403A50000E8EE432807BA00000EEC860288083A00000C;
defparam spx9_inst_6.INIT_RAM_32 = 288'h0C7074219402650000077443014402A50000067475219402E50000047443014403250000;
defparam spx9_inst_6.INIT_RAM_33 = 288'h74DE0000CCCE65000401018F1A1041E3520E186C4283ADC82009C1106E4483EDC8AB822E;
defparam spx9_inst_6.INIT_RAM_34 = 288'hF6A0101010002163D0B5A0100E175F0392E9E0705CFC0DCB9781B171F0352E1E0687FC02;
defparam spx9_inst_6.INIT_RAM_35 = 288'hC8E043280EBA000002C88602880F3A000191C48616391082C75C024C840000C042E64880;
defparam spx9_inst_6.INIT_RAM_36 = 288'h03626E219406650000016243014406A50000C4DE43280DBA000008C88602880E3A000006;
defparam spx9_inst_6.INIT_RAM_37 = 288'h0C606C219405650000076243014405A5000006626D219405E50000046243014406250000;
defparam spx9_inst_6.INIT_RAM_38 = 288'hD49E0000CACD65000401018F161041E2D20E185C4283ABC8200981105E4483EBC8AB022E;
defparam spx9_inst_6.INIT_RAM_39 = 288'h4000020B122201728040424000858A7100D9E0605AFC0BCB57817169F02D2D1E05857C02;
defparam spx9_inst_6.INIT_RAM_3A = 288'h040097248405043D51A4922A2580150E00000670131C0015614400A8F02B06000546A395;
defparam spx9_inst_6.INIT_RAM_3B = 288'h403AC600090C6622F71C002733194C45831961C858B2963CC5933965F34048060C8D8000;
defparam spx9_inst_6.INIT_RAM_3C = 288'hECF65B680000236214012EC2000EE83805B96482001B9D8EE4C0502C6800160A4542B080;
defparam spx9_inst_6.INIT_RAM_3D = 288'hD8EE4C0502C6800060281610000D9FA501D11EA03A3B1DC980A058D0000C0502C201019D;
defparam spx9_inst_6.INIT_RAM_3E = 288'hEDA00B6800006363DD401A50000086C7BE803BA000008D894F300031008BAC00003011B9;
defparam spx9_inst_6.INIT_RAM_3F = 288'h28163400030140B0804043D0080EAF6C0BD000203AA0FF000101DBEA8B1302CEE8B09DDF;

SPX9 spx9_inst_7 (
    .DO({spx9_inst_7_dout_w[26:0],spx9_inst_7_dout[17:9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[13],ad[12],ad[11]}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[17:9]})
);

defparam spx9_inst_7.READ_MODE = 1'b0;
defparam spx9_inst_7.WRITE_MODE = 2'b01;
defparam spx9_inst_7.BIT_WIDTH = 9;
defparam spx9_inst_7.BLK_SEL = 3'b011;
defparam spx9_inst_7.RESET_MODE = "SYNC";
defparam spx9_inst_7.INIT_RAM_00 = 288'hE8F00B100007009DC0ECF47D6800004363D9FBA000008D893005D7980001806DCEC77260;
defparam spx9_inst_7.INIT_RAM_01 = 288'hCBA000008C8E473280381E3000030140B0804062C90004072F9680ADA039BCD4C703FDC0;
defparam spx9_inst_7.INIT_RAM_02 = 288'h0C7277280AFA000018C8F25000401018119904013320E02744280EECF4716800004323D9;
defparam spx9_inst_7.INIT_RAM_03 = 288'h707AC00006C7AC00D8F580035D96C7AC91D11E0000008F59780517C80023AF00048DA000;
defparam spx9_inst_7.INIT_RAM_04 = 288'h2C6800080381E100800016BFDFF047AC0008F5F1373B9FF6E5AAB000200B018167078200;
defparam spx9_inst_7.INIT_RAM_05 = 288'h0F00BB25E02764009A017AC01EB07767B2B54000011B14A0092BD00003009B9D8EE4C050;
defparam spx9_inst_7.INIT_RAM_06 = 288'h7FFAC01EB150013400F5803D6002D7F9FFEB007AC8C002D7F9FFEB007ACAC300276415D9;
defparam spx9_inst_7.INIT_RAM_07 = 288'h0479880301C70000602816100800000011EB060081A100003000004D403D600F5800B5FE;
defparam spx9_inst_7.INIT_RAM_08 = 288'hE885BA3D900003CDB770001B2004D003CC58FF00FB258ECC0000201879801FE0879801FE;
defparam spx9_inst_7.INIT_RAM_09 = 288'hE8F6461D98069A05D9ECC03B2004D003CC58FF00FB3E6E8BFBB3D1047440000E8A003100;
defparam spx9_inst_7.INIT_RAM_0A = 288'h2C6800040180E10080E740BB3D980767C1D17F767A208E8D4EB000040003100E8803A21C;
defparam spx9_inst_7.INIT_RAM_0B = 288'hE000018C1F402009D90C337D00801767B3354000011B11900A2A780003009B9D8EE4C050;
defparam spx9_inst_7.INIT_RAM_0C = 288'h2C20000AF8800101DDEEA0136082079C00A4F3EC7726028163400030140B0804001004E7;
defparam spx9_inst_7.INIT_RAM_0D = 288'hE892BA3B9001CCE000E0F2556800002322740122D3000060133391CCA00E078C0000C050;
defparam spx9_inst_7.INIT_RAM_0E = 288'h41A0362000C7079237D0003BDFEECF6405D9007000018ECEC5001880063B3C1107678250;
defparam spx9_inst_7.INIT_RAM_0F = 288'h000232294017CD4000060133391CCA00E078C000100703C20100179400369B9E8F4405D1;
defparam spx9_inst_7.INIT_RAM_10 = 288'h0C40031D9E080031D9D8903B26B406C40018E0F278250E89ABA3B90076CE000E0F242680;
defparam spx9_inst_7.INIT_RAM_11 = 288'hE8F4405D1B8A2001BEFF767B202EC83B0B3800201001880063B3C14000031D9D888B8000;
defparam spx9_inst_7.INIT_RAM_12 = 288'h00766B680000236224014ECA0000601373B1DC980A058D000100703C201015F2400329B9;
defparam spx9_inst_7.INIT_RAM_13 = 288'hDEA0196082079C00A4F3F079391CCA00E078C0000C0502C20101294006003D999F664A30;
defparam spx9_inst_7.INIT_RAM_14 = 288'hECEA5001880063B3C1107678250E892BA3B10032DD00071A003001E4BB792DFE800101BD;
defparam spx9_inst_7.INIT_RAM_15 = 288'h34E80006FCC00369B1E8F4405D140B2000E1406A40018E0F27BDFEECF6405D9007000018;
defparam spx9_inst_7.INIT_RAM_16 = 288'h00063B3A911700001880063B3C100063B3A920765F280D480031C1E4F04A1D1357476200;
defparam spx9_inst_7.INIT_RAM_17 = 288'h40203DBD80065363D1E880BA3FF600037DFEECF6405D90704EE0004020031000C7678280;
defparam spx9_inst_7.INIT_RAM_18 = 288'h40707B202E880B9202E0810107340706EA30F5841017F107AC0880200C071C000200E078;
defparam spx9_inst_7.INIT_RAM_19 = 288'h301610080ECEC772602C6800040180E10080D5F47B240180E38000200C070800063C81EB;
defparam spx9_inst_7.INIT_RAM_1A = 288'h4006001D94006003D90E767DC00ECF6411D90006001D908766AB98006C77260281634000;
defparam spx9_inst_7.INIT_RAM_1B = 288'h04003B280400003001EC8003000EC878001800F640018007646DD9F1003B3D9047640000;
defparam spx9_inst_7.INIT_RAM_1C = 288'h080600187207AC04B7BC0004D60000802018F0000C0502C20100000072001D9EC823B2E7;
defparam spx9_inst_7.INIT_RAM_1D = 288'h041AC90001D240002008063C000100403000B0903D60448B8000307C00040100C7800020;
defparam spx9_inst_7.INIT_RAM_1E = 288'h000802018F000040100C0022A40F58408BB00011050001004031E0000802018004EC81EB;
defparam spx9_inst_7.INIT_RAM_1F = 288'h10040300064903D640FCA000058AC00040100C78000200806000EF207AC401F8C0009DC0;
defparam spx9_inst_7.INIT_RAM_20 = 288'hF5C035B50001B910001004031E00008020180028C81EB4074FD000313C0002008063C000;
defparam spx9_inst_7.INIT_RAM_21 = 288'hDC00040100C7800020080600057207AC01875C000F020000802018F000040100C000FA40;
defparam spx9_inst_7.INIT_RAM_22 = 288'h0008020180002C81EB004EF100048540002008063C00010040300018903D600B08800084;
defparam spx9_inst_7.INIT_RAM_23 = 288'h207AC00EF2C0014C80000802018F000040100C003CA40F58022AF000271D0001004031E0;
defparam spx9_inst_7.INIT_RAM_24 = 288'h5E6C0002008063C000100403000CC903D60064F0000B00C00040100C78000200806001BF;
defparam spx9_inst_7.INIT_RAM_25 = 288'hF000040100C0029A40F5800FA900032290001004031E0000802018005CC81EB0028E5000;
defparam spx9_inst_7.INIT_RAM_26 = 288'h80903D60218D8000E23C00040100C7800020080600127207AC0257FC001ACE0000802018;
defparam spx9_inst_7.INIT_RAM_27 = 288'h003EB50001004031E00008020180036C81EB0202D900077040002008063C000100403000;
defparam spx9_inst_7.INIT_RAM_28 = 288'h0C780002008060008F207AC21BFCC0020D40000802018F000040100C0016A40F5823CA30;
defparam spx9_inst_7.INIT_RAM_29 = 288'h0010C81EB205CCD0008D1C0002008063C00010040300034903D620CCC0001106C0004010;
defparam spx9_inst_7.INIT_RAM_2A = 288'h9C00265A0000802018F000040100C0003A40F5A029BD00049810001004031E0000802018;
defparam spx9_inst_7.INIT_RAM_2B = 288'h08063C000100403000E8903D60080A80013E9C00040100C78000200806001F7207AE0127;
defparam spx9_inst_7.INIT_RAM_2C = 288'h0C0030A40F58016B7000558D0001004031E0000802018006AC81EB0036C1000A53400020;
defparam spx9_inst_7.INIT_RAM_2D = 288'h349000170CC00040100C780002008060015F207AC008F6C002C400000802018F00004010;
defparam spx9_inst_7.INIT_RAM_2E = 288'h1004031E00008020180044C81EB0010F5000BE4C0002008063C0001004030009C903D600;
defparam spx9_inst_7.INIT_RAM_2F = 288'h0C103D7EF2C003C040000020078F59006038E000040100C001DA40F58003B10006219000;
defparam spx9_inst_7.INIT_RAM_30 = 288'h1C003BC3EECF6405D9000003044ECFA0001001763B3D11076401D12C727A3C900103D7D1;
defparam spx9_inst_7.INIT_RAM_31 = 288'hEEFFB806000023D640180E38000200C0700052F640008F58000278F59006038E00008030;
defparam spx9_inst_7.INIT_RAM_32 = 288'hF40000878F590071C00010060380050C700040774001E047AC00023C7AFB61EE000011EB;
defparam spx9_inst_7.INIT_RAM_33 = 288'hC000089D91C083B2002D3E0F1EB00023D7D91F1980008F59006038E000080380077C0004;
defparam spx9_inst_7.INIT_RAM_34 = 288'h180E38000200C0700000010005AFF7FC11EB00023D6CF7C0003C00047ADBAE0000000018;
defparam spx9_inst_7.INIT_RAM_35 = 288'h000200DEA388600080EEF7401E80D023BE8710000120006203D6000A00BBFDF0002BD440;
defparam spx9_inst_7.INIT_RAM_36 = 288'h568802018F000080301C00001FE037A80010037ABEE80ED94F90004076FB600F408021DF;
defparam spx9_inst_7.INIT_RAM_37 = 288'hF1205021640203FC014D2010079FFA60E0784022121600000000001004030004A88E6000;
defparam spx9_inst_7.INIT_RAM_38 = 288'h08120803514080703028062E000080040400501C0F0804424102814C05A9C8140A01000E;
defparam spx9_inst_7.INIT_RAM_39 = 288'hE970C084820171008040203C60024100A1F000280E07840221208140A6090400D14079E0;
defparam spx9_inst_7.INIT_RAM_3A = 288'h16108881A3F02084183F009341001702506852201010340200941804043E1E0007040042;
defparam spx9_inst_7.INIT_RAM_3B = 288'h3FA003FF0100948442117FCFC9C000480040407B4844212079441F047FCFC1E000810080;
defparam spx9_inst_7.INIT_RAM_3C = 288'h102001010408605CA534767322EF02C484020010CEC9AF090884224087FFE7E51272C49C;
defparam spx9_inst_7.INIT_RAM_3D = 288'h3F88256A04F79F448051A0081F901190848102041007C34FE4D481EB158DDED402268000;
defparam spx9_inst_7.INIT_RAM_3E = 288'h407D100800008100080820500800C21102812920101872180C7FFEBCA0101F50FD9AFE26;
defparam spx9_inst_7.INIT_RAM_3F = 288'h0136281F00B02BE01C0478015F0150006C8A0000337FE202029A02C6A01016D402021C80;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[29:0],sp_inst_8_dout[19:18]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[19:18]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b01;
defparam sp_inst_8.BIT_WIDTH = 2;
defparam sp_inst_8.BLK_SEL = 3'b000;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000021C06DF304B00030000021;
defparam sp_inst_8.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_08 = 256'hFFC0C3C3C3040CFDC050028C3C38FFFFFFFFFC2021222100000033FFFFFFFFF0;
defparam sp_inst_8.INIT_RAM_09 = 256'h3003F3CF77F77DCCC2F3CFFF70C00FFFFFFFFFFFFFFFCDA30CC3FFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_0A = 256'h3FCC43FC4C3FCF30CF10FF130F3CC33CFC30010FFC4CF7F310FCF133FCC33CFC;
defparam sp_inst_8.INIT_RAM_0B = 256'h03004FD3D3FFF03003D3FCC0C00C700C01FD3F30300134C4D30C005F4C4D30C0;
defparam sp_inst_8.INIT_RAM_0C = 256'hC0077D03003BE4FDF7DF7DF3FC0C00FBE4FF7DF7DF7CFF03003E4FF7DF7DF7FF;
defparam sp_inst_8.INIT_RAM_0D = 256'h0000C0C017F3CF7C0CC0C017FFD4711C3D33F3CD03FFCF83F3C83CFCCCCCFFC0;
defparam sp_inst_8.INIT_RAM_0E = 256'hCE0CF3DC4CCF3DC4CCF3DC4CCF3DC0CCF3DC4CCF3D4CCF3D30000C33C0F0F3FF;
defparam sp_inst_8.INIT_RAM_0F = 256'h33344CC33CD74C3FC3005C3F39E0308F033C0CF3CC33CCFC0CF033CF30CF33CC;
defparam sp_inst_8.INIT_RAM_10 = 256'h303D0C00630C130CCF3703F33C30003C30000C000C00030000C00FC4CDC300CC;
defparam sp_inst_8.INIT_RAM_11 = 256'h005FFF51C470F4CFCF340FFF3E0FCF20F3F33333FF03005FCF3DF03303003F03;
defparam sp_inst_8.INIT_RAM_12 = 256'h71333CF71333CF71333CF70333CF71333CF5333CF4C04030CF03C3CFFC000303;
defparam sp_inst_8.INIT_RAM_13 = 256'h0C0170FCFFC00F080CE780C23C0CF033CF30CF33F033C0CF3CC33CCF333833CF;
defparam sp_inst_8.INIT_RAM_14 = 256'h7CF030034F03003FFDCDFFF03004333F0330CCDF03000DCCF030000C000301F3;
defparam sp_inst_8.INIT_RAM_15 = 256'hC30C0F0C00D17345CD17347345CD17C3C3FC3010FF4F33310CCF0C00DFF03003;
defparam sp_inst_8.INIT_RAM_16 = 256'h075C307570CFC3F0C00F3CFD0300030D0D18030C358034600D180318030C30C0;
defparam sp_inst_8.INIT_RAM_17 = 256'h30C78C30FF0C004D30C0075C307570CFF075C307570CFC3F0C0075C307570CFF;
defparam sp_inst_8.INIT_RAM_18 = 256'h007C71BC300373F0C00C30CF0C00D4CC34CCD4CC34CC0CD4CCD3334CC35330C5;
defparam sp_inst_8.INIT_RAM_19 = 256'hC00D74C344CFC30030C30C8F0C003330C335D4D4CCD737F7E0CC3E3F03001B0C;
defparam sp_inst_8.INIT_RAM_1A = 256'h0C00D130F3C300CF333C3000F3D87DF187CCCF75C0C00345773FC0C000CF3DC0;
defparam sp_inst_8.INIT_RAM_1B = 256'hF301C004FFD741FDDFFD03003FC4013FF74013FF5D47CD404FFD7517FDDFFDD4;
defparam sp_inst_8.INIT_RAM_1C = 256'h703430F0C000C030CCC7FF3C330FF0C033C330C0C3007CFEC0C04FFD33013FB5;
defparam sp_inst_8.INIT_RAM_1D = 256'h00530C230CF0C00D0D0340DC340D40D7030F0C0034DC35035030F0C003435C0D;
defparam sp_inst_8.INIT_RAM_1E = 256'h0C00434F034D3DD430010D34F034F750C00330C00330C07F034F4301FC0D3D0C;
defparam sp_inst_8.INIT_RAM_1F = 256'hCF381CCCF4CF3CCD77CC0C00CDF0CE7FCCF33E7FCCF27CCCCCD030033CF5DCF4;
defparam sp_inst_8.INIT_RAM_20 = 256'h3C3000CC0CCF0C00C0CCC30C323C3001CCC733134C31CCC330CC33C300207C43;
defparam sp_inst_8.INIT_RAM_21 = 256'hC3330CC3330CC33DC30001701D030010D0C7CF0C07CC1CFC30017D30CC134C33;
defparam sp_inst_8.INIT_RAM_22 = 256'h1038CC4150380380381740E0F335840F335140F0CD4030FC0C04F0C00C3330CC;
defparam sp_inst_8.INIT_RAM_23 = 256'h3CE1F3FC00F38FADD550CFF003CF3F3FC00F3CFF003C0380C0141C1C151038D6;
defparam sp_inst_8.INIT_RAM_24 = 256'hC0C017FCC450F113C33D10CC0F10C040C3F030143D1FF003C43FC00F1410FF00;
defparam sp_inst_8.INIT_RAM_25 = 256'h10F10C0C0FC0C014FD10F10C0C0FC0C017FCC0434C04D30CF443303C4300030F;
defparam sp_inst_8.INIT_RAM_26 = 256'hD0F3FCCC30D0F3FC30CF3FC30CF3FC30C0C30F0F333300CCC00C0303F030053F;
defparam sp_inst_8.INIT_RAM_27 = 256'h003005CF3C35034C0D33C3043C10F04F003005C2F30BD0FD0C340FC0C01F0FCC;
defparam sp_inst_8.INIT_RAM_28 = 256'h3D90EC1B10CEB054346C4337D90EC0B031B10FC0C0173CE059F3833CE059F382;
defparam sp_inst_8.INIT_RAM_29 = 256'h0F90F90C28DD0E8F030050A2438543458432A0543458430A097F6430CCF397CC;
defparam sp_inst_8.INIT_RAM_2A = 256'h05404370C4370C4370F50F50C140FC0C0177CF50C14C353F030059FE3FCF3DF9;
defparam sp_inst_8.INIT_RAM_2B = 256'hCF343031170D5C71C7045C3FF00473C03004CD00C3D03005AF50C1090E43F030;
defparam sp_inst_8.INIT_RAM_2C = 256'h10F4030C30C330CC3C743C743C743C743C743C74F1D0F1D0F1D0F1D0F1D0F1D3;
defparam sp_inst_8.INIT_RAM_2D = 256'h3C643C643C643C643C643C64F190F190F190F193CF301031D70C17DF7DF7DF70;
defparam sp_inst_8.INIT_RAM_2E = 256'h78FF8FFFFFFFF1F80C73DC38150CD13F431D70C77DF7DF70F0F4030C30C330CC;
defparam sp_inst_8.INIT_RAM_2F = 256'h0C0155FC1F07C4C3DD0F743DD0FC0D03F03004375FC0C014FD0C3803E3F03001;
defparam sp_inst_8.INIT_RAM_30 = 256'h3130C33300C2CB2C3D90F4030C30F90F90FC0C01607D5F73F733F90F90C200FC;
defparam sp_inst_8.INIT_RAM_31 = 256'h303005030A005CC7B305CC7B307B30330C31333E430A03F030051F30FFFB177C;
defparam sp_inst_8.INIT_RAM_32 = 256'hC2C32C3D430403F03005FF3F3CD003CCF3FFCC4DCFCF30D3CF0D4C4DCCF03333;
defparam sp_inst_8.INIT_RAM_33 = 256'h0C080FC0C0158FF31D3D8CF310F4CF3CCF9CF50C1C0FC0C011C7D030FC0C0141;
defparam sp_inst_8.INIT_RAM_34 = 256'hDC30FFC0C01743F1310C040FC0C0144FF3133CC114CF43C433C3CC74FCCF88F5;
defparam sp_inst_8.INIT_RAM_35 = 256'h5E3FCF8CF308533D0F10CF0F3DD3F33E30CFF33374FCF310F4CF3CCF80D0FCC7;
defparam sp_inst_8.INIT_RAM_36 = 256'h4D43C0C0F033CF30434F3CF3033D3C0C05FC3005FC0C01037CCCC174C5310300;
defparam sp_inst_8.INIT_RAM_37 = 256'h000CB040300033C100C000CF0803000330200C000CC0803000330200C01433CF;
defparam sp_inst_8.INIT_RAM_38 = 256'h324000C00CC90003000324000C000EA0003000368100C000CA0403000328100C;
defparam sp_inst_8.INIT_RAM_39 = 256'h080300332C300C00CCB0C0300332C300C00CC80C03003320300C00CC80003003;
defparam sp_inst_8.INIT_RAM_3A = 256'h0C008D50403002314100C00CC50803003318200C00CC60803003318200C00CC7;
defparam sp_inst_8.INIT_RAM_3B = 256'h0CC000C0C008C7000300231C000C008C40003002310100C008C4040300239410;
defparam sp_inst_8.INIT_RAM_3C = 256'h830C430F10C0C030C0C3000870303C43FD0C0C00B0C0C0C00CF300F01F337F0F;
defparam sp_inst_8.INIT_RAM_3D = 256'h145C14400300004040C0033035C07CC30311F30C49150F0C0C0001F30C403100;
defparam sp_inst_8.INIT_RAM_3E = 256'h13047400744034052141440214540F3070355C010001400000000C0000050554;
defparam sp_inst_8.INIT_RAM_3F = 256'h1F0C33010F1CD759650415055743D73C5D1513110471D35C104100D811D14D00;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[29:0],sp_inst_9_dout[21:20]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[21:20]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b01;
defparam sp_inst_9.BIT_WIDTH = 2;
defparam sp_inst_9.BLK_SEL = 3'b000;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000000C008F304F000350011F1;
defparam sp_inst_9.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_08 = 256'hFFC0C3C3C3040CFCC1500B0C3C30FFFFFFFFFC2022222220000023FFFFFFFFF0;
defparam sp_inst_9.INIT_RAM_09 = 256'h3003F3CF77F77DCCC1F3CFFF70C00FFFFFFFFFFFFFFFCF030FC3FFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_0A = 256'h3FCC87FC8C3FCF30DF21FF230F3CC37CFC30021FFC8CF7F321FCF233FCC37CFC;
defparam sp_inst_9.INIT_RAM_0B = 256'h03004FD3D3FFF03003D3FCC0C00C700C01FD3F30300238C8E30C009F8C8E30C0;
defparam sp_inst_9.INIT_RAM_0C = 256'hC0037D03003FF4FEF3EF3EF3FC0C00FFF4FFBCFBCFBCFF03003F4FFBCFBCFBFF;
defparam sp_inst_9.INIT_RAM_0D = 256'h0000C0C017F3CF7C0CC0C017FFD8B22C3D37F3CD57FFCF8BF7C8BCFCCDCCFFC0;
defparam sp_inst_9.INIT_RAM_0E = 256'hCF0CF3DC4CCF3DC4CCF3DC4CCF3DC0CCF3DC4CCF3D8CCF3D30600C73C0F1F3FF;
defparam sp_inst_9.INIT_RAM_0F = 256'h33388CC33CE78C3FC3005C7F3DF030CF073C1CF3DC734CFC1CF073CF71CD33CC;
defparam sp_inst_9.INIT_RAM_10 = 256'h303D0C00730C030CCF7703F33C30003C30000C000C00030000C00FC8CDC300CC;
defparam sp_inst_9.INIT_RAM_11 = 256'h005FFF62C8B0F4DFCF355FFF3E2FDF22F3F33733FF03005FCF3DF03303003F03;
defparam sp_inst_9.INIT_RAM_12 = 256'h71333CF71333CF71333CF70333CF71333CF6333CF4C10031CF03C7CFFC000303;
defparam sp_inst_9.INIT_RAM_13 = 256'h0C0171FCFFC00E088CF7C0C33C1CF073CF71CD33F073C1CF3DC734CF333C33CF;
defparam sp_inst_9.INIT_RAM_14 = 256'h5CF030034F03003FFDCDFFF03005373F1330CCDF03000DCCF030000C000301F3;
defparam sp_inst_9.INIT_RAM_15 = 256'hC30C0F0C00E23388CE2338B388CE23C3C3FC3014FF4F33310CCF0C00D4F03003;
defparam sp_inst_9.INIT_RAM_16 = 256'h075C307570CFC3F0C00F3CFD0300030D0D28830C368834A20D288328831C30C0;
defparam sp_inst_9.INIT_RAM_17 = 256'h30C7CC30FF0C008E30C0075C307570CFF075C307570CFC3F0C0075C307570CFF;
defparam sp_inst_9.INIT_RAM_18 = 256'h007C713C300373F0C00C30CF0C00D4CC34CCD4CC34CC0CD4CCD3334CC35330C4;
defparam sp_inst_9.INIT_RAM_19 = 256'hC00E78C388CFC30030C30C4F0C003330C339E4E4CCE33BF3E2CC3C3F0300130C;
defparam sp_inst_9.INIT_RAM_1A = 256'h0C00E230F3C300CF333C3000F3E07DF207CCCF75C0C00389BB3FC0C000CF3DC0;
defparam sp_inst_9.INIT_RAM_1B = 256'hF381E008FFD781FE8F7D03003FC8023FF78023FF6E07CE008FFD7817FE8F7DD4;
defparam sp_inst_9.INIT_RAM_1C = 256'h703430F0C000C030CCC7FF3C330FF0C033C330C0C3007CFFC2C08FFD3B023FF6;
defparam sp_inst_9.INIT_RAM_1D = 256'h00730C030CF0C00D0D0340D0360D40D7030F0C0034DC35035030F0C003435C0D;
defparam sp_inst_9.INIT_RAM_1E = 256'h0C00534F134D3DD430014D34F134F750C00330C00330C06E134F4301B84D3D0C;
defparam sp_inst_9.INIT_RAM_1F = 256'hCF361DCCD8CF3DCD76CC0C00CDF0CF7FCCF33F7FCCF37CCCCCD030033CF5ECF4;
defparam sp_inst_9.INIT_RAM_20 = 256'h3C3000CC0CCF0C00C8CCC30C303C3001CCC733238C31CCC330CC33C300187C83;
defparam sp_inst_9.INIT_RAM_21 = 256'hC3330CC3330CD33DC3000C70CD030020E0C7CF0C07CC1CFC30027E30CC238C33;
defparam sp_inst_9.INIT_RAM_22 = 256'h1134CC6151341341341B44D0F336444D336144D0CD8030FC0C04F0C00C3330CC;
defparam sp_inst_9.INIT_RAM_23 = 256'h3851F3FC00E14F0D57504FF003853D3FC00E14FF003C0340C0141414191134D9;
defparam sp_inst_9.INIT_RAM_24 = 256'hC0C017FCD461F517C33D10CC0F10C140C3F030143E1FF003C83FC00F2820FF00;
defparam sp_inst_9.INIT_RAM_25 = 256'h10F10C100FC0C014FD10F10C100FC0C017FCD4474D45D30CF443303C4305030F;
defparam sp_inst_9.INIT_RAM_26 = 256'h00F77CCC3000F77C30CF77C30CF77C30C0C30F1F333300CCC00C0303F030053F;
defparam sp_inst_9.INIT_RAM_27 = 256'h003005CF3035134C4D3300043010C04C00300502F00BD0FD0C000FC0C01F1FCC;
defparam sp_inst_9.INIT_RAM_28 = 256'h3DD0CC1710CA3098385C4327DD0CC03031710FC0C0173CC059B3033CC059B300;
defparam sp_inst_9.INIT_RAM_29 = 256'h0FD0FD0C0C990CCF03005030C3C98385C4323098385C4303097F7430CCF397CC;
defparam sp_inst_9.INIT_RAM_2A = 256'h05303370C3370C3370FD0FD0C0C0FC0C01450FD0C0C0333F030059F43DCF39FD;
defparam sp_inst_9.INIT_RAM_2B = 256'hCF302031570C482082055C3FF00C23C03004CCC0C3D03005CFD0C0C10C33F030;
defparam sp_inst_9.INIT_RAM_2C = 256'h20F4030C30C330CC3D7434743D7434743D743474F5D0D1D0F5D0D1D0F5D0D1D3;
defparam sp_inst_9.INIT_RAM_2D = 256'h3D7434743D7434743D743474F5D0D1D0F5D0D1D3CF302031170C57EFBEFBEFB0;
defparam sp_inst_9.INIT_RAM_2E = 256'h74FF4FFFFFFFC1F40C73CC342610E53E431170C7BEFBEFB0D0F4030C30C330CC;
defparam sp_inst_9.INIT_RAM_2F = 256'h0C0155FD1F47C4C3D90F643D90F00D03F03004775FC0C015F90C3443D3F03001;
defparam sp_inst_9.INIT_RAM_30 = 256'h3030C73300C30C303D90F4030C30F90F90FC0C01747D5F62E722F90F90C340FC;
defparam sp_inst_9.INIT_RAM_31 = 256'h303005230C004CC7F304CC7F307F30330C31333E430C03F030051F30FFFC11FC;
defparam sp_inst_9.INIT_RAM_32 = 256'hC3C33C3E430C03F03005FF3F3CF007CCF3FFCC4DCFCF30D7CF0F004DCCF03333;
defparam sp_inst_9.INIT_RAM_33 = 256'h0C3C0FC0C017CFF3DC7FCCF321F5DF3CCF3CF90C3C0FC0C013C7DC30FC0C0143;
defparam sp_inst_9.INIT_RAM_34 = 256'hD830FFC0C01653BF390C3C0FC0C017CFF3F33CCF15DF47C877C7CF71FCCF3CF9;
defparam sp_inst_9.INIT_RAM_35 = 256'h5A3FCE8CF338577D1F21DF1F39C7F33CE38FF3E271FCF321F5DF3CCF3C94EF87;
defparam sp_inst_9.INIT_RAM_36 = 256'h8D47C4C1F133CF30535F3CF3133A3C0C05FC3005FC0C01037CCCC078C6310300;
defparam sp_inst_9.INIT_RAM_37 = 256'h000C90803000324200C000C90803000328200C000CA0803000328200C01433CE;
defparam sp_inst_9.INIT_RAM_38 = 256'h324200C00CE90803000364200C000C90803000324200C000C90803000324200C;
defparam sp_inst_9.INIT_RAM_39 = 256'h0403003320100C00CC80403003320100C00CC90403003324100C00CC90803003;
defparam sp_inst_9.INIT_RAM_3A = 256'h0C00CC80403003320100C00CC80403003320100C00CC80403003320100C00CC8;
defparam sp_inst_9.INIT_RAM_3B = 256'h0EC100C0C00CCB040300332C100C00CC804030033A0100C00CD8040300332010;
defparam sp_inst_9.INIT_RAM_3C = 256'hC30C430F00C0C030C0C3002C70303C83F80C0C00F0C0C0C00CF304F01F337F0F;
defparam sp_inst_9.INIT_RAM_3D = 256'h145C1500030000AC80C0033031EC7CC303B1F30EC0100F0C0C0001F30EC03B01;
defparam sp_inst_9.INIT_RAM_3E = 256'h1740300070153105000004F014540F30B0055C020001400000000C0000050554;
defparam sp_inst_9.INIT_RAM_3F = 256'h1F1C37010F1CD751550415055703D77D1D5553110431C35C104515D001C05C55;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[29:0],sp_inst_10_dout[23:22]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[23:22]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b01;
defparam sp_inst_10.BIT_WIDTH = 2;
defparam sp_inst_10.BLK_SEL = 3'b000;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000011822CB2003A2232228880;
defparam sp_inst_10.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_08 = 256'hAA80D1E1D100AEE9E002AEE81D14AAAAAAAAA81111111111111112AAAAAAAAA0;
defparam sp_inst_10.INIT_RAM_09 = 256'hA29AB82222A228A90410AAA62A808AAAAAAAAAAAAAAA8EDB658AAAAAAAAAAAAA;
defparam sp_inst_10.INIT_RAM_0A = 256'h7AA8429D453AAAA04A10A7514BAA8128AAA2910A9D45E2AA10A4B517AA8128AA;
defparam sp_inst_10.INIT_RAM_0B = 256'hAA2A1BCACAC02AA2A7CAF2AA8A9D36A8A83CACAAA291944651A8A44944651A8A;
defparam sp_inst_10.INIT_RAM_0C = 256'h8A9100AA2A7EB2B1A61A618AAAA8A9FEB2BC69869862AAAA2A7F2BC69869862A;
defparam sp_inst_10.INIT_RAM_0D = 256'hAAAAAA8A8302AB0E20AA8A83AAC66198A802A28802AEAA02828028A8E888AAAA;
defparam sp_inst_10.INIT_RAM_0E = 256'hAB8AAACA28AAACA28AAACA28AAACAA8AAACA28AAAC68AAACA221282AA200A2AA;
defparam sp_inst_10.INIT_RAM_0F = 256'hA225488A289248A8AA2A0C2AAC3881EF82AE0AAA882A28BE0AB82AAA20A8A2A8;
defparam sp_inst_10.INIT_RAM_10 = 256'h4290A8A629A4A9A6A62229A62AA2922AA292A8A4A8A4AA292A8A42D490AA2908;
defparam sp_inst_10.INIT_RAM_11 = 256'h2A0EAB198662A00A8A200ABAA80A0A00A2A3A222AAAA2A0C0AAC3882AA298790;
defparam sp_inst_10.INIT_RAM_12 = 256'h28A2AAB28A2AAB28A2AAB2AA2AAB28A2AAB1A2AAB28884A0AA88028AAAAAAAAA;
defparam sp_inst_10.INIT_RAM_13 = 256'hA8A830AABA954A0028B0E207BE0AB82AAA20A8A2F82AE0AAA882A28AA2AE2AAB;
defparam sp_inst_10.INIT_RAM_14 = 256'h08AAA2A71AAA2A7EAC8CBAAAA2A0A2AA0AA2AA8EAA2A68EAAAA292A8A4AA28A2;
defparam sp_inst_10.INIT_RAM_15 = 256'h8A088AA8A495625589562562558956A9A9AAA280AA0B2A200A8AA8A9C2AAA2A7;
defparam sp_inst_10.INIT_RAM_16 = 256'h210A92102A4A8AAA8A9E3808AA2989A44850224A91022140885022502284A088;
defparam sp_inst_10.INIT_RAM_17 = 256'h9A62E692AAA8A4651A8A610A92102A4AA210A92102A4A8AAA8A610A92102A4AA;
defparam sp_inst_10.INIT_RAM_18 = 256'hA6252A5AA29A2AAA8A6AAAAAA8A682A8A2AA82A8A2A8AA82AA8AAA2A8A0AA2A0;
defparam sp_inst_10.INIT_RAM_19 = 256'h8A492482648AAA29228A2A8AA8A9122282249090889626A680A8AA2AAA29A5A8;
defparam sp_inst_10.INIT_RAM_1A = 256'hA8A4992102AA29D0202AA2A490B8008380200800AA8A9264662AAA8A924220AA;
defparam sp_inst_10.INIT_RAM_1B = 256'h55E078047740E0095554AA2A776E011DD0E011DD1781578047740E0009555042;
defparam sp_inst_10.INIT_RAM_1C = 256'h212124AA8A6A4A92AA6227AA92A6AA8A7AA92A626A2A00776B8047748E011DD1;
defparam sp_inst_10.INIT_RAM_1D = 256'hA629A4A9A4AA8A644852148521480482125AA8A6908520120124AA8A69120848;
defparam sp_inst_10.INIT_RAM_1E = 256'hA8A6091189104002A29824411891000A8A699A8A699A8A1589152A28562454A8;
defparam sp_inst_10.INIT_RAM_1F = 256'hEAAE0898B8EAA898318AA8A9EC365F2022089B22220B2222220AA2A796701442;
defparam sp_inst_10.INIT_RAM_20 = 256'h2AA29964A64AA8A6A8A8AAAAAA2AA2986A61A91944A86A6A9AA699AA2A780169;
defparam sp_inst_10.INIT_RAM_21 = 256'h8AAAAA8AAAA80AA0AA2A4B0AB0AA291A526266A8A28A0A6AA291251964194699;
defparam sp_inst_10.INIT_RAM_22 = 256'h0868A8E008688688680E21A0AA33821A2AE021A28B80A2AAA8A1AA8A68AAAAAA;
defparam sp_inst_10.INIT_RAM_23 = 256'h28E0ABA954A38AA8400A8EA5528E2A3A954A38EA5528A9EA8A8138380E0868CE;
defparam sp_inst_10.INIT_RAM_24 = 256'hAA8A83AAB810AE0286280A8A2A0A8B828AAAA282AF8EA5528EBA954A3EBAEA55;
defparam sp_inst_10.INIT_RAM_25 = 256'h0AA0A8B82AAA8A80200AA0A8B82AAA8A83AAB8221B808618A02A28A82A2E0A2A;
defparam sp_inst_10.INIT_RAM_26 = 256'hE0A228A8A0E0A228A28A228A28A228A2828A2A0A2A2A888AA2288A22AAA2A0AA;
defparam sp_inst_10.INIT_RAM_27 = 256'h8AA2A0EAAE20891A2462E3829E0A78278AA2A0E3AB8ECAACA8B82AAA8A8B0AA9;
defparam sp_inst_10.INIT_RAM_28 = 256'hA0CAB80E0A8FE045E5382A300CAB82E0A0E0AAAA8A83AAB80C62E3AAB80C62E3;
defparam sp_inst_10.INIT_RAM_29 = 256'hAACAACA8B8CC2B8AAA2A02E383C45E5382A3E045E5382A2E0C0032A28E08C000;
defparam sp_inst_10.INIT_RAM_2A = 256'hA0E0E2E28E2E28E2E2ACAACA8B82AAA8A8308ACA8B8CAE2AAA2A0CA2288A6CAC;
defparam sp_inst_10.INIT_RAM_2B = 256'hAAA2E0A0C2A838E38E030AAAAAA8E2AAA2A10B82080AA2A0BACA8B8C2BE2AAA2;
defparam sp_inst_10.INIT_RAM_2C = 256'hE0A08A28A28A2288A830A230A830A230A830A230A0C288C2A0C288C2A0C288C2;
defparam sp_inst_10.INIT_RAM_2D = 256'hA830A230A830A230A830A230A0C288C2A0C288C2AAA2E0A0C2A8C21861861862;
defparam sp_inst_10.INIT_RAM_2E = 256'h28AA8AA2222238A8282698A811C8922B2A0C2A8061861862A0A08A28A28A2288;
defparam sp_inst_10.INIT_RAM_2F = 256'hA8A8304A068040040CA832A0CAA82A0AAAA2A1D2CAAA8A83ACA8A8CAA2AAA2A8;
defparam sp_inst_10.INIT_RAM_30 = 256'h9A9A6296224A8A2828CAA08A28A2ACAACAAAA8A82800C5159215ACAACA8A82AA;
defparam sp_inst_10.INIT_RAM_31 = 256'h9AA2A0A92A060662D920662D922D90A228A8192B2A2A0AAAA2A08B9A7AAA04AA;
defparam sp_inst_10.INIT_RAM_32 = 256'h824A24AB2A2A0AAAA2A0DAAEAAA823A8A276AA348BAAAA838AA68E14889A9A9A;
defparam sp_inst_10.INIT_RAM_33 = 256'hA8A82AAA8A828EAA8A2A8EAA10A04A298AA8ACA8A82AAA8A868148926AA8A80A;
defparam sp_inst_10.INIT_RAM_34 = 256'h48926AAA8A8202AA2CA8A82AAA8A828EAAA3AA8A004A028412828A28A98AA8AC;
defparam sp_inst_10.INIT_RAM_35 = 256'h0A3AAA8EAA2801280A104A0A28A2A62AA28EAAA228AEAA10A04A298AA880AA81;
defparam sp_inst_10.INIT_RAM_36 = 256'h8821A0886822CAAA02062CAA822A2AA8A0AAA2A0EAA8A8792AAAA32A6298AA2A;
defparam sp_inst_10.INIT_RAM_37 = 256'hA9E6A28AA2A79A8A2A8A9E6A28AA2A79A8A2A8A9E6A28AA2A79A8A2A8A8032AA;
defparam sp_inst_10.INIT_RAM_38 = 256'h928A2A8A9A6A28AA2A79A8A2A8A9E6A28AA2A79A8A2A8A9E6A28AA2A79A8A2A8;
defparam sp_inst_10.INIT_RAM_39 = 256'h28AA2A6928A2A8A9A4A28AA2A6928A2A8A9A4A28AA2A6928A2A8A9A4A28AA2A6;
defparam sp_inst_10.INIT_RAM_3A = 256'hA8A9A4A28AA2A6928A2A8A9A4A28AA2A6928A2A8A9A4A28AA2A6928A2A8A9A4A;
defparam sp_inst_10.INIT_RAM_3B = 256'hA68A226A8A9A4A28AA2A69A8A2A8A9A5A28AA2A6928A2A8A9A4A28AA2A6928A2;
defparam sp_inst_10.INIT_RAM_3C = 256'h862A09A65A6A8A42626A2A681A98916955A6A8A9AA626A8A9EAA21A04A262AA6;
defparam sp_inst_10.INIT_RAM_3D = 256'h000A02EAAA00A9A8AA8A92929C28004429A001128E0E1026A8A948B9A6829A08;
defparam sp_inst_10.INIT_RAM_3E = 256'h0305244235002440944450910002AE7A3A800EA82AA82A20A8AAA8A8AAA08000;
defparam sp_inst_10.INIT_RAM_3F = 256'h470CB3005E8EC300002280800362C33C4C000B84007493048A20404510D40900;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[29:0],sp_inst_11_dout[25:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[25:24]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b01;
defparam sp_inst_11.BIT_WIDTH = 2;
defparam sp_inst_11.BLK_SEL = 3'b000;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000020D330D3003937737640C0;
defparam sp_inst_11.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_08 = 256'h5550F9E5F9208FE8F803F4185F98000000000103000000333333315555555554;
defparam sp_inst_11.INIT_RAM_09 = 256'h62343A69001004248CA141551980C0000000000000001C27C449555555555555;
defparam sp_inst_11.INIT_RAM_0A = 256'hF061201F27306186404807C9C7861900566234821F27C21848047C9F06190056;
defparam sp_inst_11.INIT_RAM_0B = 256'h96202BCACAD569620FCAF665883F3E5880BCAD996234D25349988D0925349988;
defparam sp_inst_11.INIT_RAM_0C = 256'h8831249620FC32B410410419565883FC32BD04104106559620FF2BD041041065;
defparam sp_inst_11.INIT_RAM_0D = 256'h955565880318632E2065880318C2008084028004000C610012000050E4001565;
defparam sp_inst_11.INIT_RAM_0E = 256'h638618C200618C200618C200618C280618C200618C00618C0020280862180146;
defparam sp_inst_11.INIT_RAM_0F = 256'h844321186102218566200C018CB883EF808E02184808207E0238086120208160;
defparam sp_inst_11.INIT_RAM_10 = 256'hD0D4988D2D347D3535030D50066233066233988C988CE6233988D8F234662361;
defparam sp_inst_11.INIT_RAM_11 = 256'h200C63080202100A0010003184004800014390005596200C618CB881962367B2;
defparam sp_inst_11.INIT_RAM_12 = 256'h0801863080186308018630A01863080186300186300080A0218860051A555596;
defparam sp_inst_11.INIT_RAM_13 = 256'h98803006363FC7002032E20FBE02380861202081F808E02184808205818E1863;
defparam sp_inst_11.INIT_RAM_14 = 256'h0C19620F019620FC1C8CB559620000060000010D9620D0D1196233988CE62011;
defparam sp_inst_11.INIT_RAM_15 = 256'h1820A1988D0C043010C043043010C04D4D5662021823180006059883C219620F;
defparam sp_inst_11.INIT_RAM_16 = 256'h1102111008410859883C309496235D74E0002821D0028000A00028002845820A;
defparam sp_inst_11.INIT_RAM_17 = 256'hD35374D015988D349988D102111008418110211100841085988D102111008418;
defparam sp_inst_11.INIT_RAM_18 = 256'h8D0407566234005988D18611988D000040010000400081000100040004000010;
defparam sp_inst_11.INIT_RAM_19 = 256'h88D0220432016623461861C19883148608408202210040604001871596237598;
defparam sp_inst_11.INIT_RAM_1A = 256'h588D0C83986623F98186620D963824A382788110658834300005658836580465;
defparam sp_inst_11.INIT_RAM_1B = 256'h9EE0B8027742E09809E49620F76E009DD2E009DD0B827B8027742E029809E442;
defparam sp_inst_11.INIT_RAM_1C = 256'h3080821988DB46D213530784D1355988F84D1357662026776B802774AE009DD0;
defparam sp_inst_11.INIT_RAM_1D = 256'h8D2D347D341988D4E0C8320C832002030821988DD20C800800821988DD380C20;
defparam sp_inst_11.INIT_RAM_1E = 256'h588D0D0B0D08244262343420B0D0910988DD1988DD19880C0D09262030342498;
defparam sp_inst_11.INIT_RAM_1F = 256'hE18E008078E1848030065883ECBC7F2566599F26665B26666649620FA6B08852;
defparam sp_inst_11.INIT_RAM_20 = 256'h066237447441988D1C1C1861870662344051014D24044050D435D56620F8270D;
defparam sp_inst_11.INIT_RAM_21 = 256'h00048100048180046620C8268496234F4B5045988046005662342497444D25D1;
defparam sp_inst_11.INIT_RAM_22 = 256'h000860E000080080080C00205033800218E000220780821658835988D0004810;
defparam sp_inst_11.INIT_RAM_23 = 256'h1CE01B63FC7381C400008D8FF1CE06363FC738D8FF1C6DE5880338380E0008CE;
defparam sp_inst_11.INIT_RAM_24 = 256'h6588030638080E000C14020621020B82085962026F8D8FF1CEB63FC73EBAD8FF;
defparam sp_inst_11.INIT_RAM_25 = 256'h021020B82165880184021020B8216588030638000380003050081884082E0821;
defparam sp_inst_11.INIT_RAM_26 = 256'hE060002080E0600082060008206000820208218019198A0662A0A82859620041;
defparam sp_inst_11.INIT_RAM_27 = 256'h896200E18E000D003401E380DE037807896200E30B8DC21C20B8216588038063;
defparam sp_inst_11.INIT_RAM_28 = 256'h84C2380E020FE002C23808324C2382E080E02165880386380C01E386380C01E3;
defparam sp_inst_11.INIT_RAM_29 = 256'h21C21C20B8CC2385962002E383C02C238083E002C238082E0C2930820E9AC284;
defparam sp_inst_11.INIT_RAM_2A = 256'h00E0E0C20E0C20E0C21C21C20B8216588030C1C20B8C8E0596200C9304C10C9C;
defparam sp_inst_11.INIT_RAM_2B = 256'h4102E080C02038E38E0300855008E16562038B828A496200F1C20B8C23E05962;
defparam sp_inst_11.INIT_RAM_2C = 256'hE01088208208020084328232843282328432823210CA08CA10CA08CA10CA08C8;
defparam sp_inst_11.INIT_RAM_2D = 256'h84328232843282328432823210CA08CA10CA08C84102E080C020C24104104102;
defparam sp_inst_11.INIT_RAM_2E = 256'h380380199999B8B8201C40B800CC0307080C020104104102E010882082080200;
defparam sp_inst_11.INIT_RAM_2F = 256'h588030AE0B8240824C213084C2382E08596203D2C96588031C20B8C8E0596200;
defparam sp_inst_11.INIT_RAM_30 = 256'hD7D350D0134B8E3804C2108820821C21C21658803824C90C03001C21C20B8216;
defparam sp_inst_11.INIT_RAM_31 = 256'hD962007D2E0D0453511045351135108020841107082E085962004DD3718E00C4;
defparam sp_inst_11.INIT_RAM_32 = 256'h83483487082E08596200D18C8638010041746114C321840104478D14C056D6D6;
defparam sp_inst_11.INIT_RAM_33 = 256'h20B8216588038C18C2038E184800401405B85C20B82165880F824D965658800B;
defparam sp_inst_11.INIT_RAM_34 = 256'h4D965565880300CE1C20B8216588038C18E3860E00402002102007080405B85C;
defparam sp_inst_11.INIT_RAM_35 = 256'h0E30638E18380100800840801C201016E38C18E3080E184800401405B8C03382;
defparam sp_inst_11.INIT_RAM_36 = 256'h800101004041C18404041C18441E165880566200D65880FD2666732F63D89620;
defparam sp_inst_11.INIT_RAM_37 = 256'h83F6E289620FDB8A25883F6E289620FDB8A25883F6E289620FDB8A2588007063;
defparam sp_inst_11.INIT_RAM_38 = 256'hD38A25883F7E289620FDB8A25883F6E289620FDB8A25883F6E289620FDB8A258;
defparam sp_inst_11.INIT_RAM_39 = 256'h289620FD38A25883F4E289620FD38A25883F4E289620FD38A25883F4E289620F;
defparam sp_inst_11.INIT_RAM_3A = 256'h5883F4E289620FD38A25883F4E289620FD38A25883F4E289620FD38A25883F4E;
defparam sp_inst_11.INIT_RAM_3B = 256'h378A1365883F5E289620FD38A25883F4E289620FD38A25883F4E289620FD38A2;
defparam sp_inst_11.INIT_RAM_3C = 256'h80210D35C36588DB536620F826D4D70D70365883D35365883E180020C01D0135;
defparam sp_inst_11.INIT_RAM_3D = 256'h00080015560083F8E58836D6DCB8264E6DE0993B8E0E39B65883C4DD3781DE00;
defparam sp_inst_11.INIT_RAM_3E = 256'h030020C6300020C080003080000152F639400D00200000009455584880000000;
defparam sp_inst_11.INIT_RAM_3F = 256'h80008110FE8EC300002000000322C33C0C000B80003083008000000340C00800;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[29:0],sp_inst_12_dout[27:26]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[27:26]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b01;
defparam sp_inst_12.BIT_WIDTH = 2;
defparam sp_inst_12.BLK_SEL = 3'b000;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'h000000000000000000000000000000000000000000DD14451451728470448810;
defparam sp_inst_12.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_08 = 256'hAA97090909A32400480806E39095AAAAAAAAA91011111144444406AAAAAAAAA5;
defparam sp_inst_12.INIT_RAM_09 = 256'h8C8AB28A22A2288880A2AAAA22351AAAAAAAAAAAAAAA96D82692AAAAAAAAAAAA;
defparam sp_inst_12.INIT_RAM_0A = 256'h2A8A2294242A8A2A4A88A5090B28A928A88C88889424A0A288A48092A8A928A8;
defparam sp_inst_12.INIT_RAM_0B = 256'h28CA2140406A828CA140588A328410A3289406228C8812604923220126049232;
defparam sp_inst_12.INIT_RAM_0C = 256'h32852828CA169018A28A28A2A8A32856901628A28A28AA28CA1501628A28A28A;
defparam sp_inst_12.INIT_RAM_0D = 256'h2AAA8A3281AA8924C88A3280A24020082820228802A68A32A08328A84898AA8A;
defparam sp_inst_12.INIT_RAM_0E = 256'h8908A248288A248288A248288A248288A248288A24288A24AE0C82228CA8A2A8;
defparam sp_inst_12.INIT_RAM_0F = 256'h2AA02AA28A802A2A88CA062A24932041222488A2822208848892228A08882288;
defparam sp_inst_12.INIT_RAM_10 = 256'h2218232201848186862061A2288C84688C842321232108C842322A028888C8AA;
defparam sp_inst_12.INIT_RAM_11 = 256'hCA0289008020A0808A200A9A28CA820CA2A12262AA28CA06AA24932228C8A602;
defparam sp_inst_12.INIT_RAM_12 = 256'h20A228920A228920A228920A228920A22890A22892B832088A32A28AA0AAAA28;
defparam sp_inst_12.INIT_RAM_13 = 256'h232818A89880085308924C81048892228A0888221222488A2822208A22242289;
defparam sp_inst_12.INIT_RAM_14 = 256'h01A28CA10A28CA1AA4041AA28CA0A2A80AAAAA8628CA286AA28C84232108C8A2;
defparam sp_inst_12.INIT_RAM_15 = 256'hA26A2A2322802A00A802A02A00A802A1A1A88C82A22AA2A0688A232840A28CA1;
defparam sp_inst_12.INIT_RAM_16 = 256'h21089210225A82A2328618A828C8918428030A2A1030A00C28030A030A9626A2;
defparam sp_inst_12.INIT_RAM_17 = 256'h18604612AA232204923221089210225A221089210225A82A23221089210225A2;
defparam sp_inst_12.INIT_RAM_18 = 256'h222428588C8A2AA2322A28AA232282A8A2AA82A8A2AB2A82AA8AAA2A8A0AA6A1;
defparam sp_inst_12.INIT_RAM_19 = 256'h3228028A028A88C8A8A28A1A23285AA88AA00282AA82A2828CAA286A28C88523;
defparam sp_inst_12.INIT_RAM_1A = 256'hA32280A0AA88C84AA2A88CA21A93282132889A208A328A00226A8A32886A688A;
defparam sp_inst_12.INIT_RAM_1B = 256'hA24C934255424CA00A2828CA1544D095524D095509328934255424C2A00A2880;
defparam sp_inst_12.INIT_RAM_1C = 256'h04A0A2A23220481CA860672A1286A23232A1286448CA2A554134255424D09550;
defparam sp_inst_12.INIT_RAM_1D = 256'h2201848184A23224280A0280A02812804A2A23221280A04A04A2A232210A0128;
defparam sp_inst_12.INIT_RAM_1E = 256'hA3220108810828808C8804208810A2023221923221923200810A08C802042823;
defparam sp_inst_12.INIT_RAM_1F = 256'h4A24C808934A28081088A3284492450A88A2210888A1088888828CA3289088A0;
defparam sp_inst_12.INIT_RAM_20 = 256'h288C8864864A2322A1A1A28A28688C886A61A98124A86A6A1A861988CA132821;
defparam sp_inst_12.INIT_RAM_21 = 256'h9AAA2A8AAA2A8AA888CA13283828C8804862662322880A688C88049864812619;
defparam sp_inst_12.INIT_RAM_22 = 256'hC823884C082382382346208CAA113208E24C208C893228A8A320A23228AAA2AA;
defparam sp_inst_12.INIT_RAM_23 = 256'h214CA18800853A18410A36200214E8D8800853620021814A3280131344C82344;
defparam sp_inst_12.INIT_RAM_24 = 256'h8A3280A89308A4C292284888CA48813492A28C80810620021418800854106200;
defparam sp_inst_12.INIT_RAM_25 = 256'h48A488138A8A3282A848A488138A8A3280A8932209308248A12223292204D24A;
defparam sp_inst_12.INIT_RAM_26 = 256'h4C822B8B204C822A2C8822A2C8822A2C88A28A8A222232888C8A22CAA28CA0AA;
defparam sp_inst_12.INIT_RAM_27 = 256'h328CA04A24E0810A04224D3214C85325328CA04DA13648A488138A8A32898A88;
defparam sp_inst_12.INIT_RAM_28 = 256'h28489344C8854C00201322128489304E244C8A8A3281289304224D289304224D;
defparam sp_inst_12.INIT_RAM_29 = 256'h8A48A4881344093A28CA004D3140020132214C0020132204C42A122C8CA2428B;
defparam sp_inst_12.INIT_RAM_2A = 256'hA04C4E6C84E6C84E6CA48A488130A8A328101A48813424EA28CA0420681A2424;
defparam sp_inst_12.INIT_RAM_2B = 256'hAAA04E244288134D34D10A2AAAA34E8A8CA0813CB2828CA05A488134094EA28C;
defparam sp_inst_12.INIT_RAM_2C = 256'h4CA0328A28B2288A281220122812201228122012A0488048A0488048A048804A;
defparam sp_inst_12.INIT_RAM_2D = 256'h281220122812201228122012A0488048A048804AAAA04E244288408A28A28A20;
defparam sp_inst_12.INIT_RAM_2E = 256'h13A93AAAAAAA901388228813000180692244288228A28A204CA0328A28B2288A;
defparam sp_inst_12.INIT_RAM_2F = 256'hA32810A4C9328082848A1228489304E2A28CA050428A3281A48813424EA28CA8;
defparam sp_inst_12.INIT_RAM_30 = 256'h18186212244134D32848A0124A28A48A48A8A32813284A008040A48A488138A8;
defparam sp_inst_12.INIT_RAM_31 = 256'h128CA08104C2166059216605920592228A2859692204E2A28CA081185A24C02A;
defparam sp_inst_12.INIT_RAM_32 = 256'h317217292204E2A28CA09A262893A1A8A2668A14198A2A818A95361418981818;
defparam sp_inst_12.INIT_RAM_33 = 256'h88138A8A32813AA248293CA288A04A288A13A488138A8A328132861868A32801;
defparam sp_inst_12.INIT_RAM_34 = 256'h86186A8A32810664E488138A8A32813AA24F2884C04A22A212A28920A88A13A4;
defparam sp_inst_12.INIT_RAM_35 = 256'h04EA893CA21301288A884A8A2482A2284D3AA24D20ACA288A04A288A13419932;
defparam sp_inst_12.INIT_RAM_36 = 256'h3821A1A868629A2A060629A28624E8A320A88CA068A3281108888504411028CA;
defparam sp_inst_12.INIT_RAM_37 = 256'h28444C328CA11130CA328444C328CA11130CA328444C328CA11130CA32836689;
defparam sp_inst_12.INIT_RAM_38 = 256'h1530CA328444C328CA11130CA328444C328CA11130CA328444C328CA11130CA3;
defparam sp_inst_12.INIT_RAM_39 = 256'hC328CA11530CA328454C328CA11530CA328454C328CA11530CA328454C328CA1;
defparam sp_inst_12.INIT_RAM_3A = 256'hA328454C328CA11530CA328454C328CA11530CA328454C328CA11530CA328454;
defparam sp_inst_12.INIT_RAM_3B = 256'h8530E44A328454C328CA11530CA328454C328CA11530CA328454C328CA11530C;
defparam sp_inst_12.INIT_RAM_3C = 256'h328A1186084A32286448CA13281918218084A32868644A328CA2E08C0A222A86;
defparam sp_inst_12.INIT_RAM_3D = 256'h420242EAA80328534A32881814932A42814CA90934040A84A3280811853214F8;
defparam sp_inst_12.INIT_RAM_3E = 256'h0100020410000010000001004202A408729002A9CAA82A6129AAA3A32AA08400;
defparam sp_inst_12.INIT_RAM_3F = 256'h018611900000000410C280904008002000000000110004030A20004044400000;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[29:0],sp_inst_13_dout[29:28]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[29:28]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b01;
defparam sp_inst_13.BIT_WIDTH = 2;
defparam sp_inst_13.BLK_SEL = 3'b000;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000110041040524450448814;
defparam sp_inst_13.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_08 = 256'hAA90094909602440480406609090AAAAAAAAA95055555500000002AAAAAAAAA4;
defparam sp_inst_13.INIT_RAM_09 = 256'h808AA28A22A2288880A6AAAA22000AAAAAAAAAAAAAAA96482782AAAAAAAAAAAA;
defparam sp_inst_13.INIT_RAM_0A = 256'h2A8A2290246A8A2A4A88A4091A28A929A88088889024A0A288A58092A8A929A8;
defparam sp_inst_13.INIT_RAM_0B = 256'h280A2140406A8280A140588A028010A028940622808812604920220126049202;
defparam sp_inst_13.INIT_RAM_0C = 256'h028528280A169018A28A28A2A8A02856901628A28A28AA280A1501628A28A28A;
defparam sp_inst_13.INIT_RAM_0D = 256'h2AAA8A0280AA8924498A0282A240240A28602A9802A28A12A08129A948A8AA8A;
defparam sp_inst_13.INIT_RAM_0E = 256'h8918A248298A248298A248298A248298A248298A24298A24A204822284A8A6A8;
defparam sp_inst_13.INIT_RAM_0F = 256'h2AA02AA28A802A2A880A022A24912446222888A28222099888A2228A08882689;
defparam sp_inst_13.INIT_RAM_10 = 256'h2218202201858186862061A228808028808020202020080802022A02888808AA;
defparam sp_inst_13.INIT_RAM_11 = 256'h0A0A89009028A180AA600A8A284A8204A6A522A2AA280A02AA2491262808A502;
defparam sp_inst_13.INIT_RAM_12 = 256'h20A628920A628920A628920A628920A62890A628928812088A12A29AA0AAAA28;
defparam sp_inst_13.INIT_RAM_13 = 256'h202808A888801841089244911888A2228A0888266222888A2822209A26246289;
defparam sp_inst_13.INIT_RAM_14 = 256'h01A280A10A280A1AA4141AA280A0A2A84AAAAA86280A286AA2808020200808A2;
defparam sp_inst_13.INIT_RAM_15 = 256'hA22A2A2022802A00A802A02A00A802A1A1A88082A229A2A4289A202840A280A1;
defparam sp_inst_13.INIT_RAM_16 = 256'h61089610224AA2A2028658A82808918428010A2A1010A00428010A010A9622A2;
defparam sp_inst_13.INIT_RAM_17 = 256'h18604612AA202204920221089610224A261089610224AA2A20221089610224A2;
defparam sp_inst_13.INIT_RAM_18 = 256'h22242858808A2AA2022A28AA202282A9A2AA82A9A2A92A82AA8AAA2A9A0AA2A1;
defparam sp_inst_13.INIT_RAM_19 = 256'h0228029A028A8808A8A28A1A20285AA88AA00282AA82A28284AA286A28088520;
defparam sp_inst_13.INIT_RAM_1A = 256'hA02280A0AA88080AA6A880A21A91282512889A208A028A00226A8A02886A688A;
defparam sp_inst_13.INIT_RAM_1B = 256'hA2449182554244A00A28280A15446095524609550912891825542442A00A2880;
defparam sp_inst_13.INIT_RAM_1C = 256'h04A0A2A202205814A860652A1686A20212A16864480A2A554118255424609550;
defparam sp_inst_13.INIT_RAM_1D = 256'h2201858184A20224280A0280A02812804A2A20221280A04A04A2A202210A0128;
defparam sp_inst_13.INIT_RAM_1E = 256'hA022010881082880808804208810A2020221920221920200810A080802042820;
defparam sp_inst_13.INIT_RAM_1F = 256'h8A244809918A28081098A0284482450A88A2210888A10888888280A2289089A0;
defparam sp_inst_13.INIT_RAM_20 = 256'h28808865864A2022A1A1A28A286880886A61A98124A86A6A1A8619880A112821;
defparam sp_inst_13.INIT_RAM_21 = 256'hAAAA2AAAAA2A8AA8880A1128182808804862662022980A688088049865812619;
defparam sp_inst_13.INIT_RAM_22 = 256'h482189440821821821062085AA41120862442084991524A8A020A2022AAAA2AA;
defparam sp_inst_13.INIT_RAM_23 = 256'h6144A08801851A18410A122006146848801851220061814A0280515104482104;
defparam sp_inst_13.INIT_RAM_24 = 256'h8A0282A89108A442826848984A489118A2A28080850220061408801854102200;
defparam sp_inst_13.INIT_RAM_25 = 256'h48A489114A8A0282A848A489114A8A0282A8912209108209A12261292244628A;
defparam sp_inst_13.INIT_RAM_26 = 256'h45822A8A2545822A289822A289822A2894924A8A626212988489224AA280A0AA;
defparam sp_inst_13.INIT_RAM_27 = 256'h1280A08A2460810A04264512144851251280A045A11648A489114A8A02888A88;
defparam sp_inst_13.INIT_RAM_28 = 256'h2848910448954400201122528489144520448A8A028228910426462891042645;
defparam sp_inst_13.INIT_RAM_29 = 256'h8A48A4891144891A280A0445154002011225440020112244542A122498A24299;
defparam sp_inst_13.INIT_RAM_2A = 256'hA04546649466494664A48A489118A8A028101A489116246A280A0420681A2424;
defparam sp_inst_13.INIT_RAM_2B = 256'hAAA445204289114514410A2AAAA1468A80A09118A28280A05A4891148946A280;
defparam sp_inst_13.INIT_RAM_2C = 256'h44A1228A2892288A281220122812201228122012A0488048A0488048A048804A;
defparam sp_inst_13.INIT_RAM_2D = 256'h281220122812201228122012A0488048A048804AAAA445204289408A28A28A24;
defparam sp_inst_13.INIT_RAM_2E = 256'h11A91AAAAAAA901149228911000180692204289228A28A2444A1228A2892288A;
defparam sp_inst_13.INIT_RAM_2F = 256'hA02810A449128082848A122848914452A280A050428A0281A489116246A280A8;
defparam sp_inst_13.INIT_RAM_30 = 256'h18186212645114512848A1228A28A48A48A8A02811284A008040A48A489114A8;
defparam sp_inst_13.INIT_RAM_31 = 256'h1280A0814452166059616605960595224A285929224452A280A081184A24402A;
defparam sp_inst_13.INIT_RAM_32 = 256'h15525529224452A280A09A2A289161A9A6668A141A8A2A819A95161419981818;
defparam sp_inst_13.INIT_RAM_33 = 256'h89114A8A02811AA2482918A288A04A689A11A489114A8A028112861868A02811;
defparam sp_inst_13.INIT_RAM_34 = 256'h86186A8A028106646489114A8A02811AA2462894404A229212A29920A89A11A4;
defparam sp_inst_13.INIT_RAM_35 = 256'h046A8918A25101288A484A8A6482A268451AA24520A8A288A04A689A11419912;
defparam sp_inst_13.INIT_RAM_36 = 256'h1821A19868669A2A060669A2866468A020A880A068A02811088885044110280A;
defparam sp_inst_13.INIT_RAM_37 = 256'h2844441280A111104A02844441280A111104A02844441280A111104A02806689;
defparam sp_inst_13.INIT_RAM_38 = 256'h15104A02844441280A111104A02844441280A111104A02844441280A111104A0;
defparam sp_inst_13.INIT_RAM_39 = 256'h41280A115104A02845441280A115104A02845441280A115104A02845441280A1;
defparam sp_inst_13.INIT_RAM_3A = 256'hA02845441280A115104A02845441280A115104A02845441280A115104A028454;
defparam sp_inst_13.INIT_RAM_3B = 256'h8510644A02845441280A115104A02845441280A115104A02845441280A115104;
defparam sp_inst_13.INIT_RAM_3C = 256'h128A1186084A022864480A11281918218084A02868644A0288A220840A622A86;
defparam sp_inst_13.INIT_RAM_3D = 256'h4102426AA80028514A02881814912A428144A90914040A84A028181185161448;
defparam sp_inst_13.INIT_RAM_3E = 256'h8200011400008010000001008102A418529006A90AA82A2128AAA1A02AA0A400;
defparam sp_inst_13.INIT_RAM_3F = 256'h0186115004044104100280904104422404000000500000000A20004040000000;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[29:0],sp_inst_14_dout[31:30]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:30]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b01;
defparam sp_inst_14.BIT_WIDTH = 2;
defparam sp_inst_14.BLK_SEL = 3'b000;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000004500000000104010000004;
defparam sp_inst_14.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_08 = 256'h0001404040410440400400010400000000000054555555444444400000000000;
defparam sp_inst_14.INIT_RAM_09 = 256'h0400100000000000100400000010000000000000000004010000000000000000;
defparam sp_inst_14.INIT_RAM_0A = 256'h1000000400500000000001001100000100040000040040000001100100000100;
defparam sp_inst_14.INIT_RAM_0B = 256'h0040014040400004014050001004100100140400040000000001000000000010;
defparam sp_inst_14.INIT_RAM_0C = 256'h1004000040141010000000000001005410140000000000004015014000000000;
defparam sp_inst_14.INIT_RAM_0D = 256'h0000001001000104410010010040040100400410000400100001010140110000;
defparam sp_inst_14.INIT_RAM_0E = 256'h0110004001000400100040010004001000400100040100040400400004000400;
defparam sp_inst_14.INIT_RAM_0F = 256'h0000000000000000004004000411044500040000000001140010000000000401;
defparam sp_inst_14.INIT_RAM_10 = 256'h0000010000010000000000004004000004000100010000400010004000004000;
defparam sp_inst_14.INIT_RAM_11 = 256'h4004010010040100104000100040000404050044000040040004110400400100;
defparam sp_inst_14.INIT_RAM_12 = 256'h0004001000400100040010004001000400100400101001000010001000000000;
defparam sp_inst_14.INIT_RAM_13 = 256'h0100100010001011011044111400100000000004500040000000001004044001;
defparam sp_inst_14.INIT_RAM_14 = 256'h0000040100004014041410000400000040040004004000400004000100004000;
defparam sp_inst_14.INIT_RAM_15 = 256'h0041000100000000000000000000000000000400000100044010010040000401;
defparam sp_inst_14.INIT_RAM_16 = 256'h4000040000101000100451000040000000010000001000040001000100000410;
defparam sp_inst_14.INIT_RAM_17 = 256'h0000000400010000001000000400001004000040000101000100000040000100;
defparam sp_inst_14.INIT_RAM_18 = 256'h0000000004000000100000000100000100000001000100000000000010000400;
defparam sp_inst_14.INIT_RAM_19 = 256'h1000001000100040000000000100400010000000000000000400000000400001;
defparam sp_inst_14.INIT_RAM_1A = 256'h0100000400004040040004000010000500011000001000000040001000004000;
defparam sp_inst_14.INIT_RAM_1B = 256'h0040104011004000000000401104100440410044010001040110040000000000;
defparam sp_inst_14.INIT_RAM_1C = 256'h0000000010001004000001000400001010004000004000110104011004100440;
defparam sp_inst_14.INIT_RAM_1D = 256'h0000010001001000000000000000000000000100000000000000001000000000;
defparam sp_inst_14.INIT_RAM_1E = 256'h0100000000000000040000000000000010000010000010000000004000000001;
defparam sp_inst_14.INIT_RAM_1F = 256'h4004000110400000101001004410050000000100000100000000040100100100;
defparam sp_inst_14.INIT_RAM_20 = 256'h4004000100100100000000000000040000000000010000000000000040100000;
defparam sp_inst_14.INIT_RAM_21 = 256'h1000001000000000004010000000400000000001001040000400000001000000;
defparam sp_inst_14.INIT_RAM_22 = 256'h0000014000000000004400010051000000400000110504000100001001000000;
defparam sp_inst_14.INIT_RAM_23 = 256'h4040010001010000410004000404001000101040004000401000505044000044;
defparam sp_inst_14.INIT_RAM_24 = 256'h0010010010000400104040104040110410000400050400040410001014104000;
defparam sp_inst_14.INIT_RAM_25 = 256'h4004011040001000004004011040001001001000010000410100410100441040;
defparam sp_inst_14.INIT_RAM_26 = 256'h4100010105410001041000104100010414104000404010100401004000040000;
defparam sp_inst_14.INIT_RAM_27 = 256'h0004004004000000000441000400100100040041010440040110400010010000;
defparam sp_inst_14.INIT_RAM_28 = 256'h0040104400154100001000500401044104400000100100100404410010040441;
defparam sp_inst_14.INIT_RAM_29 = 256'h0040040110444100004004410550000100054100001000441400100414004011;
defparam sp_inst_14.INIT_RAM_2A = 256'h0041404414044140440400401104000100100040110504000040040000000404;
defparam sp_inst_14.INIT_RAM_2B = 256'h0004410440011041041100000000400004001104100004005040110441400004;
defparam sp_inst_14.INIT_RAM_2C = 256'h4101104104104411001000100010001000100010004000400040004000400040;
defparam sp_inst_14.INIT_RAM_2D = 256'h0010001000100010001000100040004000400040000441044001400000000004;
defparam sp_inst_14.INIT_RAM_2E = 256'h1001000000001010410001104000000100440010000000044101104104104411;
defparam sp_inst_14.INIT_RAM_2F = 256'h0100100401000000040010004010441000040040400010010401105040000400;
defparam sp_inst_14.INIT_RAM_30 = 256'h0000000040110410404001104104040040000100100040000000040040110400;
defparam sp_inst_14.INIT_RAM_31 = 256'h0004000044100000004000000400050441000041004410000400000010040000;
defparam sp_inst_14.INIT_RAM_32 = 256'h0510510100441000040040040010400104100000010000001001040001000000;
defparam sp_inst_14.INIT_RAM_33 = 256'h0110400010010400400104000000004010100401104000100100040000010011;
defparam sp_inst_14.INIT_RAM_34 = 256'h0400000010010044040110400010010400410014000000100000110000101004;
defparam sp_inst_14.INIT_RAM_35 = 256'h0410010400500000004000004400004041040041000400000000401010401100;
defparam sp_inst_14.INIT_RAM_36 = 256'h0000001000044000000044000044000100000400400100100000010401000040;
defparam sp_inst_14.INIT_RAM_37 = 256'h0040400004010100001004040000401010000100404000040101000010011001;
defparam sp_inst_14.INIT_RAM_38 = 256'h0100001004040000401010000100404000040101000010040400004010100001;
defparam sp_inst_14.INIT_RAM_39 = 256'h0000401010000100404000040101000010040400004010100001004040000401;
defparam sp_inst_14.INIT_RAM_3A = 256'h0100404000040101000010040400004010100001004040000401010000100404;
defparam sp_inst_14.INIT_RAM_3B = 256'h0100000010040400004010100001004040000401010000100404000040101000;
defparam sp_inst_14.INIT_RAM_3C = 256'h0040000000001000000040100000000000000100400000100400400100400000;
defparam sp_inst_14.INIT_RAM_3D = 256'h4100400000010050401000000410001000400041044440000100100001040410;
defparam sp_inst_14.INIT_RAM_3E = 256'h4110011010004000001000044100001050100401400000450100000100001401;
defparam sp_inst_14.INIT_RAM_3F = 256'h0041004404044104104000104104411404000100411005010000000004400000;

SP sp_inst_15 (
    .DO({sp_inst_15_dout_w[27:0],sp_inst_15_dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[13],ad[12]}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]})
);

defparam sp_inst_15.READ_MODE = 1'b0;
defparam sp_inst_15.WRITE_MODE = 2'b01;
defparam sp_inst_15.BIT_WIDTH = 4;
defparam sp_inst_15.BLK_SEL = 3'b010;
defparam sp_inst_15.RESET_MODE = "SYNC";
defparam sp_inst_15.INIT_RAM_00 = 256'h20CFF4C4DE4EF4EE0E04E4EDEF00804D3C7581FCD0DC0004004C0FFC04C5DCD5;
defparam sp_inst_15.INIT_RAM_01 = 256'hD000EF0FF0054DDDDCE4ECCCC0C50C4F4CDDC0C5F44DD4EDDCDC5540FDCDE0DD;
defparam sp_inst_15.INIT_RAM_02 = 256'hF0FF0E0E0FF4E44DCCC0EC050CFF4C4DE4EF4EE0E04E4EDEF00054DDDD0C0CEE;
defparam sp_inst_15.INIT_RAM_03 = 256'hCD0DDDCEECFC05F44ECCF4EEF0FF0E0E0F51FC4D4CE4E04EEFEF4E4F000E0E0F;
defparam sp_inst_15.INIT_RAM_04 = 256'h0F0C15CFE0E2F24FF5CFCC540F00F0CEC4E0E00EFF000054DEDD0DC054DDD0DC;
defparam sp_inst_15.INIT_RAM_05 = 256'hF5F44554CDCDDDFC1EECECE00F5FC4D4CE4E04EEFEF4E4ECE00F0FCEEDF5CE4E;
defparam sp_inst_15.INIT_RAM_06 = 256'h0C1CEECF1CFCEEC0F5C1EECF5F5CF3C40F44D44E4EEEFF000E0E0F44D44E4EEE;
defparam sp_inst_15.INIT_RAM_07 = 256'h33E0EEEFCE4EFC1EECF1FFC40EFFE4F12FC40FEC1C000FCE4DF5CE4E0F5F3C4F;
defparam sp_inst_15.INIT_RAM_08 = 256'hEEEF0C1CFEFCE04FDFC5EECFCEEC0F5FCCFCF3C4F0CCEECF51FFC4FCE04DF44C;
defparam sp_inst_15.INIT_RAM_09 = 256'hEE22207EF4D0C1FDF1DD05FE000FC0EFCEFECDCDFFFFC4FCEEDCDCDEF44C33E0;
defparam sp_inst_15.INIT_RAM_0A = 256'hFFECC4CEFD41CC0C20D434DDDDDD4C15054DDDDCEF3F4ED0020DDFFD3F420E2F;
defparam sp_inst_15.INIT_RAM_0B = 256'h0D1CF42D0F40DC010F4D000C1E20DE00E01F4002EE4F34204F020054DCDDFDE3;
defparam sp_inst_15.INIT_RAM_0C = 256'h014441ED41244D170470465EE1CD0F1173FFCE3E054DDDDF3EEEF4ED0F40DCF4;
defparam sp_inst_15.INIT_RAM_0D = 256'h9EFD9DFD70F970CD4DCD4FF44F47F4F44B44BAF4D87974140F1AEDFAFDF70DA7;
defparam sp_inst_15.INIT_RAM_0E = 256'hEFD41CC0C20D4CCDDEF4DDDDFFF8F865FFD58945DFCC4F6ED464D4709670FDDC;
defparam sp_inst_15.INIT_RAM_0F = 256'hC0DC0CD0EDEEEDEDEDFFC0ECFCEF10D0CEEC0DC00CC0FE0D003547DDDDFECC4C;
defparam sp_inst_15.INIT_RAM_10 = 256'h0F1F12CDDEEDF12D0FFD0FCFDF420F1DFD4D44C4FC1DFDCDF2E3E3230FEDECFE;
defparam sp_inst_15.INIT_RAM_11 = 256'hC0DC00CC0FEDC0FC0F8D24CE2FFF0FCFCEFDEDD0C4D20F12DCDEEDFD144C04F4;
defparam sp_inst_15.INIT_RAM_12 = 256'h007060D40DD7251E0FDCFEDECFEC0DC0CD0EDEEEDEFFFC8FFC0ECFCEF10D0CEE;
defparam sp_inst_15.INIT_RAM_13 = 256'hCEEE05CD00F271F75C7F7CC070FE0F77C4CFF6F047CC004704757470D4006C0D;
defparam sp_inst_15.INIT_RAM_14 = 256'hFD04054DDDD4CEDDDDDD14C30F6DE02F00EE00E4306F2DF0DD00007DF1E24CEC;
defparam sp_inst_15.INIT_RAM_15 = 256'h2ECF12E4F6DE0054D4DDEDCF12EC04F622FDD4034F0400FF71DE2F2C4CFD0FE0;
defparam sp_inst_15.INIT_RAM_16 = 256'h14C50044EC8849C56C0E9C6987DA9B9EF74713FE3CCD054DDDDE4C3CF3F6EFF1;
defparam sp_inst_15.INIT_RAM_17 = 256'hFF41CEEBE1FE77CC900EDE05E11CC76454B445BBCE8DF61E164F81166E05EE88;
defparam sp_inst_15.INIT_RAM_18 = 256'hCDD0D4C4DFFD0DEE0354987DDDDEC44DEDECDD0D4C4DFFD0DEEC44E4D0DCEE99;
defparam sp_inst_15.INIT_RAM_19 = 256'hFDDDFDFDFE4DC4F4CE0DFCEEEC0FEDDE4DE40FFF4CECE4EFFD3D3F3FEC44DEDE;
defparam sp_inst_15.INIT_RAM_1A = 256'hF4CEF4CEFDFECCDFE4DC4F4CE0DFCEEEC0FEDDE4DE40FFF4FEFECFC4D4CE4F0D;
defparam sp_inst_15.INIT_RAM_1B = 256'hEF2CFCDFCC4C4FCF12C04747192785E3102CDECE00FEFECFC4D4CE4F0DFDDDFD;
defparam sp_inst_15.INIT_RAM_1C = 256'h2C04054DDDDEFFCDEEF0FE0ECDCEFFE0E3DCCEEC0EED0DE3CFFE0EF0EED0EDDC;
defparam sp_inst_15.INIT_RAM_1D = 256'h0054DDDD0EEFFC000FC0CC0704CFDCECCEDEE0FE030EDDCEC29C9FCDD4C4CDC1;
defparam sp_inst_15.INIT_RAM_1E = 256'hF410C0CF3DDC2CEDCDFCDD4C4CDC4DD0C0C054F0EFEFC0C00C0C00770F410C0C;
defparam sp_inst_15.INIT_RAM_1F = 256'h0FEFFCFCFDFF0FFDED3D054DFDD0DE054DDD0DEED0CCC4EFFCFE03DC9CDED9CC;
defparam sp_inst_15.INIT_RAM_20 = 256'hCEECD0D000FEFFCCECDF3DDC2CEDCDFCDD4C4CDCCECD04FEFFCF0E5EFF0FDDFC;
defparam sp_inst_15.INIT_RAM_21 = 256'hEFDFECECD0FDC0FEFCFF3F3ED8EC0FCC29CDCDDDF4DD0C0C0FFC29C0C000F3DC;
defparam sp_inst_15.INIT_RAM_22 = 256'hE8DCDCCCF5D9EC0FDDFC0FEFCFF5DDECF5EFFC000FEFFCF3D8ECF0E5FECFF5EF;
defparam sp_inst_15.INIT_RAM_23 = 256'hCFFE5EFFFCCE8DCDCCCF5EFFFEFFCF3DEEFED8EC0F0EFEFCF3D9ECFEFF0D0FCC;
defparam sp_inst_15.INIT_RAM_24 = 256'h88888888C6273057000004CC04544E4CCFE0FEEFDE0400444CEC5DECFE0FFD9E;
defparam sp_inst_15.INIT_RAM_25 = 256'h888888888C4C8888888888888888888888888888888888888888CCCCCCCCC488;
defparam sp_inst_15.INIT_RAM_26 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC0000000008CCCCCCCCCC048848888448;
defparam sp_inst_15.INIT_RAM_27 = 256'h5D527DD1DD080408455DD5202D020465D8CC8CCCC88CCCCCCCCCC080CCCCCCCC;
defparam sp_inst_15.INIT_RAM_28 = 256'hDDE2CB404B05809BD6A090902D09C3D198094090DF5D7CD0D7DA952200A80434;
defparam sp_inst_15.INIT_RAM_29 = 256'hC055B083B840DB640204D562CBD50204D562CBD34D0EF0B08F34DDDE2CB4934D;
defparam sp_inst_15.INIT_RAM_2A = 256'h13D270482B0993D17270487B09C53DD120B0940B740B04D45B57051B94D4D5BD;
defparam sp_inst_15.INIT_RAM_2B = 256'h49B0F73FB334FB034FB033FB134FB9394B45004D9BDF3DC93FB030C4B523DDB1;
defparam sp_inst_15.INIT_RAM_2C = 256'h84CCC08CC088C880C048C40CCC04CCC4C8C4C8C4C8C4844C84C0C88408C0CB0E;
defparam sp_inst_15.INIT_RAM_2D = 256'h03DA0880C48CC448CCC4C8C0C4CCC0C8CC44C880084CC48CCC84C44048404088;
defparam sp_inst_15.INIT_RAM_2E = 256'h01A8090AAE2C01A80A5A0D04001A000DDEDDC30301DAA3001AA4D5502A59AA49;
defparam sp_inst_15.INIT_RAM_2F = 256'h00809F48003480044AEAA040060204006D5E101AE5E79E5E8790562C01A0562C;
defparam sp_inst_15.INIT_RAM_30 = 256'h045A445A04035A03095A87095A096A001200190000500001000A8080DB020048;
defparam sp_inst_15.INIT_RAM_31 = 256'h05A3D0E1240D83009C840AE0F0000EEC4FE0F000F49847A250A03E05A000E387;
defparam sp_inst_15.INIT_RAM_32 = 256'hC404DD2052FD30BA3DA3E4307DD3DDD5DC03A55CCA3D524A3D52E124FD30F4EF;
defparam sp_inst_15.INIT_RAM_33 = 256'h02255604A60530FDD0C9A42B30530024E3549804044F3A4D0405003D0D9040E4;
defparam sp_inst_15.INIT_RAM_34 = 256'h9EC53DA004DA4249201A8D15171727048701A57A3D0A1E437D40C8DDDD24A505;
defparam sp_inst_15.INIT_RAM_35 = 256'hA8DD01901AF03E2D0FDF007C30C401A41CD0CA6DD4028169C2803060F9C30CDE;
defparam sp_inst_15.INIT_RAM_36 = 256'h3D410DA45DA455DEDFD4320431A02C101A5484023AA41AE1101AAE439A02C901;
defparam sp_inst_15.INIT_RAM_37 = 256'h83150429524100DEEE3EEEAAEEE94EEEAA0E3A84AAEEEE6EEEA00555E0D0C8F0;
defparam sp_inst_15.INIT_RAM_38 = 256'h58CCCCCCCCCCCCCCCC048C048C048C048C048C048C048C048CA050C503083050;
defparam sp_inst_15.INIT_RAM_39 = 256'h89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF;
defparam sp_inst_15.INIT_RAM_3A = 256'hFF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C;
defparam sp_inst_15.INIT_RAM_3B = 256'h5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89FF5C89;
defparam sp_inst_15.INIT_RAM_3C = 256'h000000000000000C4C00010849030888000000000448000000880404048803C8;
defparam sp_inst_15.INIT_RAM_3D = 256'h00000000000000000000000000000000000BC4E0100000000000000000000000;
defparam sp_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_16 (
    .DO({sp_inst_16_dout_w[27:0],sp_inst_16_dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[13],ad[12]}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]})
);

defparam sp_inst_16.READ_MODE = 1'b0;
defparam sp_inst_16.WRITE_MODE = 2'b01;
defparam sp_inst_16.BIT_WIDTH = 4;
defparam sp_inst_16.BLK_SEL = 3'b010;
defparam sp_inst_16.RESET_MODE = "SYNC";
defparam sp_inst_16.INIT_RAM_00 = 256'hF8E86688A0888AC0D0D00AAA00E12BDE98EAEBC8A9EA002002800F9028A8A088;
defparam sp_inst_16.INIT_RAM_01 = 256'h8CEAA8EEA02AC20808C88E8EAB0A8E8E888088800A0A088A0A0AAA09C80C84A4;
defparam sp_inst_16.INIT_RAM_02 = 256'hFD00C0CA0F8C8A88E8EB001A8EE8888A0888AC0D0D00AAA00E12AC2080B808C8;
defparam sp_inst_16.INIT_RAM_03 = 256'h80ACA0EC8E98008C88888600FD00C0CA0FE1A88A8808678C0C0C008CF1CEC8AE;
defparam sp_inst_16.INIT_RAM_04 = 256'h0FB8100D8C45696F9A808EA81491FB8C888CACA8F0B002AC20081002AC208108;
defparam sp_inst_16.INIT_RAM_05 = 256'hF00800AA8A8800FA1CCAE8010FE888A8808678C0C0C008E801AE0F8C88F08C88;
defparam sp_inst_16.INIT_RAM_06 = 256'hB81ACCAD10FA8CACFEA18CAF090E89860F80AD8C08A0FCF1CEC80F80AD8C08A0;
defparam sp_inst_16.INIT_RAM_07 = 256'hD7CF680F8C88FA18CAF188A8CEE866F198A80F081ECE0F8888F088880F08786F;
defparam sp_inst_16.INIT_RAM_08 = 256'h680FB810D8F88A88AFAECCAFACCA0F0E8E9E8986FB8ACCAF0188A8F88C88F808;
defparam sp_inst_16.INIT_RAM_09 = 256'hCCDF1EEEE00D8F20E9C0CAAA000F010F8CE88E808F8886F8CC88C808F808D7CF;
defparam sp_inst_16.INIT_RAM_0A = 256'hF8282A0000038E829A80B080808084DE2A86EC0000BF10A41DAAAE6EB01D1C1E;
defparam sp_inst_16.INIT_RAM_0B = 256'h10F8F1DA0F01002F0F0011509C1DC8EDE2FF11F1C47415DCFC4D02A860EC000B;
defparam sp_inst_16.INIT_RAM_0C = 256'hA99989889959F8D0AB0AACC2C50218DD76F00C1E2A86EC00BC20F10A0F0100F0;
defparam sp_inst_16.INIT_RAM_0D = 256'hAA8AAAE80AAC0AAC0A8A9AA99889E489966F2E80E49243980E3EE2EEEAE0A8C0;
defparam sp_inst_16.INIT_RAM_0E = 256'h000038E829A808E8888D8CEAEA0EE0EEE0EAEA9E88889E88E989290AAC0AAAA8;
defparam sp_inst_16.INIT_RAM_0F = 256'h09201C81CA820C0C0AF001AA3000B9A90800820110838080026A876EC08282A0;
defparam sp_inst_16.INIT_RAM_10 = 256'h0FBF398A8A08F99C0F180F8E22990F9EAC2A8889F8B8EAC0FD6DC7F10F800090;
defparam sp_inst_16.INIT_RAM_11 = 256'h08201108380001FE0F48F984F4FA0FEF000C0A0800010F39A88A08FA388809FA;
defparam sp_inst_16.INIT_RAM_12 = 256'h080C0C8E8C8EDA9EFA0AF80009009201C81CA820C0F9FE4F001AA3000B9A9080;
defparam sp_inst_16.INIT_RAM_13 = 256'h88A0AAAA00F305F8EA0FA80F0F080F88E0CFD0D2EE8002E02EE8A0AA8E8C0CAE;
defparam sp_inst_16.INIT_RAM_14 = 256'hA8892A86C80100202020DFAF0F00CE5A0CCC1504B10C5A0FACBF1EEEE10B9808;
defparam sp_inst_16.INIT_RAM_15 = 256'h100F1109F00C02A861C8000F110089F0550CE6F1ECA0BEAFE1E05E181C0C1C88;
defparam sp_inst_16.INIT_RAM_16 = 256'h398A19192210598888BC322970AA887EEF9796F0B8802A86C800181EFBF0CCF1;
defparam sp_inst_16.INIT_RAM_17 = 256'hE29320C2EFAC9F8E4D9C8CBC23908FC9A1A9BA6C4CD2CC3AFCD28D3C26BA0C0C;
defparam sp_inst_16.INIT_RAM_18 = 256'h8AEA8B8B8A08A80826A87776C80C8B98A088AEA8B8B8A08A80889B898A8CCCE2;
defparam sp_inst_16.INIT_RAM_19 = 256'hE888A0A0F0BAEF1100FCECA80AC8AA808888CE0F9C88CB0FC6DA701FC8B98A08;
defparam sp_inst_16.INIT_RAM_1A = 256'hF100F100A0F0880F0BAEF1100FCECA80AC8AA808888CE0F4F800A90B8180B81A;
defparam sp_inst_16.INIT_RAM_1B = 256'hCE50E2248090900475001A7E1C5E8AAB1FD88CEA00F800A90B8180B81AE888A0;
defparam sp_inst_16.INIT_RAM_1C = 256'h50012AEA0C0AEA8ACECD06CACAC8C08C81EC0CE89C001CCD08E01E8ACAACAC00;
defparam sp_inst_16.INIT_RAM_1D = 256'h02AEA0C09CC88CE864C8868A874FACAC88ACE70017CAA88C8508224A090B0047;
defparam sp_inst_16.INIT_RAM_1E = 256'hF998884F142258C0800CA090B00C980888C6E1F9CEC8C8486C8078AE0F998884;
defparam sp_inst_16.INIT_RAM_1F = 256'h0FCE8CF8EA800FDE8A7E2AEA00C1002AEA0C10CC08E807A8A8D801A82ACC2000;
defparam sp_inst_16.INIT_RAM_20 = 256'h0EC081A9F1F48C40C00F1A8858C0800CA090B00C0C0061FCE8CF9C00F8EAAC00;
defparam sp_inst_16.INIT_RAM_21 = 256'hCEACCAC0E88C48F4E4CF1D1AC8C00F805A2A8240F980888C0F8050218351F108;
defparam sp_inst_16.INIT_RAM_22 = 256'hC80880C0FEC242EAAC000F4E4CFEC242FE48C4E80FC88CF1C0C0F9CEE44CF00F;
defparam sp_inst_16.INIT_RAM_23 = 256'h0F0C0EF8F80C80880C0F00F8F48C4F1ACEDAC8C00F9C84C4F1C242FCE8EC0F80;
defparam sp_inst_16.INIT_RAM_24 = 256'h00000000E66330770000288E28C8088A80A1EC00A02002A8EC0CAA0AF010FC8C;
defparam sp_inst_16.INIT_RAM_25 = 256'h0000000000A70000000000000000000000000000000000000000888888888000;
defparam sp_inst_16.INIT_RAM_26 = 256'h33333333333333333333333333333333CCCCCCCCC333333333332B00D0700B40;
defparam sp_inst_16.INIT_RAM_27 = 256'h602750262207262766600272700336760E3303A33E733333333334DB33333333;
defparam sp_inst_16.INIT_RAM_28 = 256'h2567356075067274250000006000670303303303047076000700027522073664;
defparam sp_inst_16.INIT_RAM_29 = 256'h6066506656702576272626773566272626773567620667506676625673567766;
defparam sp_inst_16.INIT_RAM_2A = 256'h6627626675066626776266750666625677506725772506576577066576576656;
defparam sp_inst_16.INIT_RAM_2B = 256'h7650567557765507755077556775567675770272756565667550603656662556;
defparam sp_inst_16.INIT_RAM_2C = 256'h8796C615C5F4C303C201C07FCE7ECDBDCC3CA9997606547321E1FEDEED4D4504;
defparam sp_inst_16.INIT_RAM_2D = 256'h076000B0CFDFCFAECDBDCCBCCB8ACA29C828C7776504C3E2C17100D0FDFDCAE9;
defparam sp_inst_16.INIT_RAM_2E = 256'h2607203006732607232006262260000036036727040006726006666250200060;
defparam sp_inst_16.INIT_RAM_2F = 256'h2232665322753227536002722527272250736260266662666660677326006773;
defparam sp_inst_16.INIT_RAM_30 = 256'h2670547006057007047067267006700266023322233222332220327355052276;
defparam sp_inst_16.INIT_RAM_31 = 256'h7637002677706622066720626222236376626222566676074700725700706667;
defparam sp_inst_16.INIT_RAM_32 = 256'h6626006267606263700627725607060706233763637067737027267760625736;
defparam sp_inst_16.INIT_RAM_33 = 256'h3336762673266260676607766067227766676426077673662606227626726027;
defparam sp_inst_16.INIT_RAM_34 = 256'h6336400326006766726073626767762667260663700362776022112222363222;
defparam sp_inst_16.INIT_RAM_35 = 256'h0730236260626276760423424336260666022370662723522523355252243603;
defparam sp_inst_16.INIT_RAM_36 = 256'h6076700660077606660777777600736260267727600760366260027760073626;
defparam sp_inst_16.INIT_RAM_37 = 256'h7637077667567502224222002224522200364367002224422200227262002762;
defparam sp_inst_16.INIT_RAM_38 = 256'h62555555555555550572D84FA51C72E94FB61C83E950B62D8307626624076370;
defparam sp_inst_16.INIT_RAM_39 = 256'h6665666665666665666665666665666665666665666665666665666665666665;
defparam sp_inst_16.INIT_RAM_3A = 256'h6566666566666566666566666566666566666566666566666566666566666566;
defparam sp_inst_16.INIT_RAM_3B = 256'h6666656666656666656666656666656666656666656666656666656666656666;
defparam sp_inst_16.INIT_RAM_3C = 256'h000009000000000D700020C11C045111AB2BA2BBAAA639998655806080570766;
defparam sp_inst_16.INIT_RAM_3D = 256'h000000000000000000000000000000000000E300000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_17 (
    .DO({sp_inst_17_dout_w[27:0],sp_inst_17_dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[13],ad[12]}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11:8]})
);

defparam sp_inst_17.READ_MODE = 1'b0;
defparam sp_inst_17.WRITE_MODE = 2'b01;
defparam sp_inst_17.BIT_WIDTH = 4;
defparam sp_inst_17.BLK_SEL = 3'b010;
defparam sp_inst_17.RESET_MODE = "SYNC";
defparam sp_inst_17.INIT_RAM_00 = 256'h19DD225818CA29105C50014DC0C8ACC5C100CC44DD000000001803C801555C45;
defparam sp_inst_17.INIT_RAM_01 = 256'h51501D194A011E210D1C51DF8CC4DD111050C1C02109640101C4510C19C14A16;
defparam sp_inst_17.INIT_RAM_02 = 256'hF16C9ED10F51D1441DFC00C45D1CC5818CA29101C50010DC08C011E210C10D50;
defparam sp_inst_17.INIT_RAM_03 = 256'h50114CD1C59C02514DD5C22C31EC5ED10F0112218D80AE9D0DC500D1DC5D9DC4;
defparam sp_inst_17.INIT_RAM_04 = 256'h03C1000189EE252B14C2DF94E604FC11D0511DCD5A420011E021C00011E21C01;
defparam sp_inst_17.INIT_RAM_05 = 256'h70040641011460FD110581C003050018D80AE9D09C500DC1C0C40BD50572D105;
defparam sp_inst_17.INIT_RAM_06 = 256'hC11D105100FD905DF1D19057894DDC52074011212A90F1DCDD1D034011212A90;
defparam sp_inst_17.INIT_RAM_07 = 256'hD211A9C3D1057D190531D21EDD9522F1D21E03CD0F510BD40572D8050F4D252B;
defparam sp_inst_17.INIT_RAM_08 = 256'hA9CBC1005CFDC50513D11053D1050B41DFDDDC52FC1D105741D21EFD4905B0CD;
defparam sp_inst_17.INIT_RAM_09 = 256'h94D9C9C00005C5E0D4DC9C00000F0C03DD155550CBD052FD51555504F0CDD211;
defparam sp_inst_17.INIT_RAM_0A = 256'hBCE96D00C822DF52D9D00EC44C082210011E11000C0B80926911D109CC0CE905;
defparam sp_inst_17.INIT_RAM_0B = 256'hC010FC0D078C00E10700A4E0410514D5521B0E1082E2064155E90011E0110000;
defparam sp_inst_17.INIT_RAM_0C = 256'h866A8AECAE2612008508511A1202E1D5003CCD0F011E110C01A0F405074000BC;
defparam sp_inst_17.INIT_RAM_0D = 256'h9DD9DD1208500851E11D191E2C2CEDE0E114122292E2224009A59E9151108640;
defparam sp_inst_17.INIT_RAM_0E = 256'h0C822DF52D5D4516EAD164555D211115514411AC11D1A9E2DAE612085C085599;
defparam sp_inst_17.INIT_RAM_0F = 256'hE5202554519AA1C501302ED5A004D111250E16E2E09A5A44000110E110CE9650;
defparam sp_inst_17.INIT_RAM_10 = 256'h0B136D15150D30950B9A03D16E59070959E1899DF0D41114B8AC92140B900E50;
defparam sp_inst_17.INIT_RAM_11 = 256'hE16E2E09A5A4C4F1076A1A9A96F1031B00090148CC40076D51190DB1A8990D31;
defparam sp_inst_17.INIT_RAM_12 = 256'hCC00A94195DC0C0000C03100ED0E5202554519AA9CF4B16B02ED52004D111250;
defparam sp_inst_17.INIT_RAM_13 = 256'h4D5C5C0000360E3544C705C501210FDC4CDB8A1000DC000800444C014110ADD1;
defparam sp_inst_17.INIT_RAM_14 = 256'h5521012E110000E4AC280110038091E901112066CC0C2D0514D1CDC00005C909;
defparam sp_inst_17.INIT_RAM_15 = 256'h000FCC00F4050012E011C00F8C00617062041E105416599DC000604001210545;
defparam sp_inst_17.INIT_RAM_16 = 256'hA2202212E6221511991933EE021111021120203C0150012E110CCD0F707CD0B4;
defparam sp_inst_17.INIT_RAM_17 = 256'h5D66EADE9D8CDEDE511151012A135606C0C64C10D115C4EDE11D6420ED08999D;
defparam sp_inst_17.INIT_RAM_18 = 256'h5DF51111250E1E0C0012000E110DD1E55805DF51111250E1E0C5A1D669115555;
defparam sp_inst_17.INIT_RAM_19 = 256'h16585C50B01DD52004D115150D1DD9481E2859470181D14BC6CD2247DD1E5D80;
defparam sp_inst_17.INIT_RAM_1A = 256'hB00CB000503C150701DD5E004D115150D1DD9481E2899432FD00DA0D209ADE4D;
defparam sp_inst_17.INIT_RAM_1B = 256'h9120511210DC5C06A2028824AC2CCC90C04D4D0000B900D60D209ADE4D16581C;
defparam sp_inst_17.INIT_RAM_1C = 256'h2028011C210D15D9DF5DC65D111150D1D0510199550AC5D10D12C1511511D51D;
defparam sp_inst_17.INIT_RAM_1D = 256'h0011C210E1DD05D566119668566F51D1559DFE00C6DD9119524D516109C50066;
defparam sp_inst_17.INIT_RAM_1E = 256'hB121E16F2611A514D51510DC50011EC9ED160EFE11D05961E1DA62040B1A5E56;
defparam sp_inst_17.INIT_RAM_1F = 256'h07D105F959D80315DDAF011C021C00011C21C015099AC2DD5D1D02555D59156C;
defparam sp_inst_17.INIT_RAM_20 = 256'h09565611143ED0625C032955A514D515101C5001E5C06E3D1053E100D5DDD915;
defparam sp_inst_17.INIT_RAM_21 = 256'hD5151510510561BE160F894D11950F9421112560716C1E910B94221221207009;
defparam sp_inst_17.INIT_RAM_22 = 256'h155521103051A1DDD9150FE1607051A1B0ED06510FDD05B411957E101E60D007;
defparam sp_inst_17.INIT_RAM_23 = 256'h57CD0FB079015552110B00D53ED06B49DFDD11950BE1DE063451A13D50D50B90;
defparam sp_inst_17.INIT_RAM_24 = 256'hFFFFFFFFD03840010000011E045481C1569C11CC9000000CF141C080B0C07559;
defparam sp_inst_17.INIT_RAM_25 = 256'hFFFFFFFFFDCDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEFF;
defparam sp_inst_17.INIT_RAM_26 = 256'h77777777777777777777777777777777666666666677777777776DFFCFCFFDDF;
defparam sp_inst_17.INIT_RAM_27 = 256'h1A8D1AD3ED05D1C52F6AA0011A088453A5775747755777777777754577777777;
defparam sp_inst_17.INIT_RAM_28 = 256'hD05E1410D5080005D13050506A0505A119709309A6EAE9A0AEA058D1A1008455;
defparam sp_inst_17.INIT_RAM_29 = 256'h1032400840F0D6007519DE1E1D402519DE1E1D140D04D08052340D05E1444340;
defparam sp_inst_17.INIT_RAM_2A = 256'h40DE1C49090240DE4E1C490902530D0C50902D474D4201055701039405055035;
defparam sp_inst_17.INIT_RAM_2B = 256'h0D509086386D23005730055330D9340405090C4DD309F01E8630F0E52410D014;
defparam sp_inst_17.INIT_RAM_2C = 256'hAAEA9AEA9A6A9A6A9A5A9A499939990999E999B999B99949999988888848DE05;
defparam sp_inst_17.INIT_RAM_2D = 256'h0A13CC8C9BCB9BCB9B9B9B7B9B6B9B9B9B6B9B5BBBDB9B3B9B2BBB0BAAFAAAEA;
defparam sp_inst_17.INIT_RAM_2E = 256'hD7005080D5E1470059000EC2C470000A05A05DD402A4DD087001D065F9359DA0;
defparam sp_inst_17.INIT_RAM_2F = 256'h0080DC38003380023A34055140A4351400D04670A251CA2551C0E1E1D700E1E1;
defparam sp_inst_17.INIT_RAM_30 = 256'hCF308F300F0330030E30EECE300E1305C101000006000020000080080505302E;
defparam sp_inst_17.INIT_RAM_31 = 256'h5401A0E2095AF840AC0F0003500000E3870450094F40F55E250080F300F058EE;
defparam sp_inst_17.INIT_RAM_32 = 256'h1941AA5E01EAEC501A0A1E4515A0A3A3AECAD3AD101A30901A47E2092AECD104;
defparam sp_inst_17.INIT_RAM_33 = 256'h240D3FD1D830C25A019E051080E303050910EAD10E003D0DD10E430D8D9D1009;
defparam sp_inst_17.INIT_RAM_34 = 256'hD04C0A0201A04520C9700048D4E4E1C4909703001A052E140A444469384A5000;
defparam sp_inst_17.INIT_RAM_35 = 256'h0D0AAF457025F0051EA17C00F0E5270043A400AA318569810F469C28910F9AA0;
defparam sp_inst_17.INIT_RAM_36 = 256'hFA1D9A0F3A0143A507AA412A4300E13370840122B3014004437000A4400E1437;
defparam sp_inst_17.INIT_RAM_37 = 256'h56010E2E109C850EEEEEEEEDEEECFEEEE0858B9FDDEEE44EEEE0E3E450A05C25;
defparam sp_inst_17.INIT_RAM_38 = 256'h8AAAAAAAAAAAAAAAAA77666555544433322221110000FFFEEE0429524F056010;
defparam sp_inst_17.INIT_RAM_39 = 256'h1227851227851227851217851217851217851217851217851217851217851217;
defparam sp_inst_17.INIT_RAM_3A = 256'h3785123785123785123785123785123785122785122785122785122785122785;
defparam sp_inst_17.INIT_RAM_3B = 256'h8512478512478512478512478512478512478512478512478512378512378512;
defparam sp_inst_17.INIT_RAM_3C = 256'h00000C00000000033300004004006666446446444446CAAAACAAABCBABAC0151;
defparam sp_inst_17.INIT_RAM_3D = 256'h000000000000000000000000000000000000E230000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_18 (
    .DO({sp_inst_18_dout_w[27:0],sp_inst_18_dout[15:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[13],ad[12]}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:12]})
);

defparam sp_inst_18.READ_MODE = 1'b0;
defparam sp_inst_18.WRITE_MODE = 2'b01;
defparam sp_inst_18.BIT_WIDTH = 4;
defparam sp_inst_18.BLK_SEL = 3'b010;
defparam sp_inst_18.RESET_MODE = "SYNC";
defparam sp_inst_18.INIT_RAM_00 = 256'h8DD39133CB33C3484739E573F044A18384DDFFFF8888000000000FC0001910B9;
defparam sp_inst_18.INIT_RAM_01 = 256'hF9E654EF020007500818FBFF8FF04D0191113210B19333B389701803E77618E1;
defparam sp_inst_18.INIT_RAM_02 = 256'hA04F1F150881F108BFF000F03D3C433CB33C348F739E5D3F0410007500F80838;
defparam sp_inst_18.INIT_RAM_03 = 256'h31932F838F9100818F33C58FB03FFF95070039133BB43B338A739E409F1F9491;
defparam sp_inst_18.INIT_RAM_04 = 256'h02F8000249D39351B31BFF8333C38F8188FF5D544F0E00007050F00000750F08;
defparam sp_inst_18.INIT_RAM_05 = 256'hD0019983B3833328038F74F00003D533BB43B3389739E444F0F10C838FD0818F;
defparam sp_inst_18.INIT_RAM_06 = 256'hF80838F3001838FF208038F1030D4C35013DC1918334F04F0F740C3DC1918334;
defparam sp_inst_18.INIT_RAM_07 = 256'h4C483331818F28038FB039343D339570393409FF016C0A838FB0838F0D049351;
defparam sp_inst_18.INIT_RAM_08 = 256'h3332F800F318398F538038F5838F040BFF5D4C35BF8838FB003934C8308F53CB;
defparam sp_inst_18.INIT_RAM_09 = 256'h4F84F4F8D00083308F0FCF8D00020F07838F3FBE333D35A838F3FBE363CB4C48;
defparam sp_inst_18.INIT_RAM_0A = 256'h6F84F700FF0BFF1E81190F5090C00000000750000F0C000A0100BB0593083400;
defparam sp_inst_18.INIT_RAM_0B = 256'hF3002000000F2021020033903875E1BD191A0C403EC8751ED1E1000070500000;
defparam sp_inst_18.INIT_RAM_0C = 256'h0143F11F31A3CC10090018C3AE00F0013CDFFF010007500F0831E0000C0010D0;
defparam sp_inst_18.INIT_RAM_0D = 256'h88F313CC00930019F3D35BC2C5C3B3B538C221202818CC4C03FCCF323C800940;
defparam sp_inst_18.INIT_RAM_0E = 256'h0FF0BFF1E8518008D0F503391302C8CA1C322213C83C3F45F313C8009300123F;
defparam sp_inst_18.INIT_RAM_0F = 256'h13CB13B83833F874E1B0388FC000D04C11132B133B33B7700040037500F84F10;
defparam sp_inst_18.INIT_RAM_10 = 256'h040D3810FE13E0BC0F110FF58F8F020894F13C44433B34E7243C45E7086013A0;
defparam sp_inst_18.INIT_RAM_11 = 256'h32B133B33B70F0E0011103F3C8B00809000EE106FE00093801FA1381F3C407F0;
defparam sp_inst_18.INIT_RAM_12 = 256'h24031301832F0F0D88FD860139013CB13B83833F7771605D0388FF000D04C111;
defparam sp_inst_18.INIT_RAM_13 = 256'hF89F0F8D00D70E8110F939FA032C0B110F1BB1C0039F000000110F5301131531;
defparam sp_inst_18.INIT_RAM_14 = 256'hD1010007500000F000F000000C0008F1000CA000930843004F85F1F8D0008303;
defparam sp_inst_18.INIT_RAM_15 = 256'h01020F30700000007050F0070F2051D03403EB8751DD181EF0803D330E387514;
defparam sp_inst_18.INIT_RAM_16 = 256'h2CB46C53538C56CC93518C33208CC8158C83CCDF08310007500FFF0190400010;
defparam sp_inst_18.INIT_RAM_17 = 256'h314AD32AB2355B3124C4BAC423C332C1DDA6A25C28C3B4322C8344B313C33911;
defparam sp_inst_18.INIT_RAM_18 = 256'hBFF1E05D111321AF04001237500F858F7F0BFF1E05D1113211F835F082E3A22B;
defparam sp_inst_18.INIT_RAM_19 = 256'h833F87EEF0588F1000D03B11132B133B1B17730C53B53E7333C31E7BF858F9F0;
defparam sp_inst_18.INIT_RAM_1A = 256'h900FA0002E6F831D0588FE000D03B11132B133B1B17830F086013A013DB33B83;
defparam sp_inst_18.INIT_RAM_1B = 256'h43DB33D358373BE27305F440F83F8F3DFDF8F88800530137013DB33B83833F57;
defparam sp_inst_18.INIT_RAM_1C = 256'h30F3000750083F8BFFDFF09D03B1113210B3B433B388704703EA761BE182D3B3;
defparam sp_inst_18.INIT_RAM_1D = 256'h00007500F8838FE4A225F0C8802E83F308BFF600F0DD3A242DA33D358473BE23;
defparam sp_inst_18.INIT_RAM_1E = 256'h004AF02203B333DB33D358373BE203FAF324047F8388F12082CF02800A032FE2;
defparam sp_inst_18.INIT_RAM_1F = 256'h05838F5333B307CB1F3F0007050F00000750F0831B38F083F85100828F34A28F;
defparam sp_inst_18.INIT_RAM_20 = 256'hBB83B384438838FD3F0A04A233DB33D358473BE233F0F41838FBF800F36D34B2;
defparam sp_inst_18.INIT_RAM_21 = 256'h838F3FBE328F2D883F8B080D2A420B4AD3B38335004FBF420C4AD3B384452003;
defparam sp_inst_18.INIT_RAM_22 = 256'hD3B38335A02B32DD34B20A83F8803B32D0838F8B0F838FC02B42BF8038F8C005;
defparam sp_inst_18.INIT_RAM_23 = 256'h26FF01F8C3AD3B3833570083B838FA0BFFBD2A4208F8388FD02B323838CF0C3A;
defparam sp_inst_18.INIT_RAM_24 = 256'h1111111110633376000000BF019131B3B1B7334C3200001FF272F8FDB0F092A4;
defparam sp_inst_18.INIT_RAM_25 = 256'h1111111111111111111111111111111111111111111111111111111111111111;
defparam sp_inst_18.INIT_RAM_26 = 256'h2222222222222222222222222222222222222222222222222222211111111111;
defparam sp_inst_18.INIT_RAM_27 = 256'h6073602662023622757003266007766602222222222222222222222222222222;
defparam sp_inst_18.INIT_RAM_28 = 256'h2073663056070376264020205002060330330330056066000600273606227666;
defparam sp_inst_18.INIT_RAM_29 = 256'h6077707670602700766623636630666623636637220662606776720736637767;
defparam sp_inst_18.INIT_RAM_2A = 256'h6223636626037223636366260367220662603577657706067776077606066266;
defparam sp_inst_18.INIT_RAM_2B = 256'h0560676676657707677076677756777727060362560660666670606667602066;
defparam sp_inst_18.INIT_RAM_2C = 256'hAA5AAA5AAA5AAA5AAA5AAA5AAA5AAA5AAA4AAA4AAA4AAA4AAA4AAA4AAA4A5405;
defparam sp_inst_18.INIT_RAM_2D = 256'h0366AA4AAA6AAA6AAA6AAA6AAA6AAA6AAA6AAA6AAA6AAA6AAA6AAA6AAA5AAA5A;
defparam sp_inst_18.INIT_RAM_2E = 256'h6622203307366622203203373662000027026037040206266202626740720032;
defparam sp_inst_18.INIT_RAM_2F = 256'h2273665732657327507506666507766650626762077660776660363666203636;
defparam sp_inst_18.INIT_RAM_30 = 256'h3662666206066206066236366206660266033222332223322222732722064276;
defparam sp_inst_18.INIT_RAM_31 = 256'h6726002726606672062622277222226667267220767266527720606620606636;
defparam sp_inst_18.INIT_RAM_32 = 256'h6676006626603362600362756600070703336736626062626066272670336626;
defparam sp_inst_18.INIT_RAM_33 = 256'h3630762603326670066606626026772627726726022276262602772662726026;
defparam sp_inst_18.INIT_RAM_34 = 256'h62662003360066773662036736363636626626226002726720BBBB6676632303;
defparam sp_inst_18.INIT_RAM_35 = 256'h2030027762766006660342525266662076062230662632232435225244252300;
defparam sp_inst_18.INIT_RAM_36 = 256'h6066700660067606260076707720367762762677660662266762020772036776;
defparam sp_inst_18.INIT_RAM_37 = 256'h2726027662666602222222202224522220766446202225522220376662002276;
defparam sp_inst_18.INIT_RAM_38 = 256'h7777777777777777777777777777777777777777777766666607766756027260;
defparam sp_inst_18.INIT_RAM_39 = 256'h6766766766766766766766766766766766766766766766766766766766766766;
defparam sp_inst_18.INIT_RAM_3A = 256'h6676676676676676676676676676676676676676676676676676676676676676;
defparam sp_inst_18.INIT_RAM_3B = 256'h7667667667667667667667667667667667667667667667667667667667667667;
defparam sp_inst_18.INIT_RAM_3C = 256'h00000B0000000001110010A11A00999999999999999988888888888888880766;
defparam sp_inst_18.INIT_RAM_3D = 256'h000000000000000000000000000000000000D130000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_19 (
    .DO({sp_inst_19_dout_w[27:0],sp_inst_19_dout[19:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[13],ad[12]}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[19:16]})
);

defparam sp_inst_19.READ_MODE = 1'b0;
defparam sp_inst_19.WRITE_MODE = 2'b01;
defparam sp_inst_19.BIT_WIDTH = 4;
defparam sp_inst_19.BLK_SEL = 3'b010;
defparam sp_inst_19.RESET_MODE = "SYNC";
defparam sp_inst_19.INIT_RAM_00 = 256'h627121157257771050020545F121110505EE44440033000500500FF005533034;
defparam sp_inst_19.INIT_RAM_01 = 256'h0545552F01055FE3565404FE2FF02750200000057525777104001357F30003F0;
defparam sp_inst_19.INIT_RAM_02 = 256'hD54F4F250E4505044FEF55F017020057257771030020525F112055FE35F3045C;
defparam sp_inst_19.INIT_RAM_03 = 256'h5055EF4540D005454000200FE54F2F350D55121157257771040020554F5F3521;
defparam sp_inst_19.INIT_RAM_04 = 256'h0DF3555C5271211FC104FEC75771DF354C035325FF000055F5E3F55055FE3F53;
defparam sp_inst_19.INIT_RAM_05 = 256'hD55527F5330571E455C0D5F10D5020057257771030020535F1010E45C0E545C0;
defparam sp_inst_19.INIT_RAM_06 = 256'hF3545C0B55D45C01D5455C0C0D0702000C5275330571E52F3F250A5275330571;
defparam sp_inst_19.INIT_RAM_07 = 256'h5330571C45C0C455C09512111711219512110CFF50000C45C0C545C00901211B;
defparam sp_inst_19.INIT_RAM_08 = 256'h5719F355A5B450C05B455C0B45C00B04FEB702009F345C08051211B451C0B527;
defparam sp_inst_19.INIT_RAM_09 = 256'h5400F143E5500551042F143E00085F5A45C0544F5D0200A45C0544F5C5275330;
defparam sp_inst_19.INIT_RAM_0A = 256'hFF650F55FF04FD0846045F0010F05555055FE3555F5F05010500470250501510;
defparam sp_inst_19.INIT_RAM_0B = 256'hF055E0500E0F05050E5510457000F04F005E5F057F400004F0050055F5E35555;
defparam sp_inst_19.INIT_RAM_0C = 256'h0110F44F000540CA01A01F450455F5440FFFFF50055FE35F5350D0500D0505D0;
defparam sp_inst_19.INIT_RAM_0D = 256'h33F00504A01CA013F1211220004533200F4CC0C01FCF445000F33F0050FA01CA;
defparam sp_inst_19.INIT_RAM_0E = 256'h5FF04FD08420305323F0205330000F4204C0CC1C4F500F33F0050FA01CA0110F;
defparam sp_inst_19.INIT_RAM_0F = 256'h0572153F30570F0B01A55460A55075020000070552777000000550FE35F65005;
defparam sp_inst_19.INIT_RAM_10 = 256'h0C590400F900C5FF0DEE0B05404B0D5000F0020DB75771F0B75771F00FF500F5;
defparam sp_inst_19.INIT_RAM_11 = 256'h007055277700F0F50DDD50F020C50C5D55500100FF050D0400FD00C0F0200FB5;
defparam sp_inst_19.INIT_RAM_12 = 256'h005050050004545E33FEFF500F50572153F30570F0FFF5FC55460C5507502000;
defparam sp_inst_19.INIT_RAM_13 = 256'h401F143E00FF5FF530FF53FF500F0F530F0FF5F0553F005005530F0005005005;
defparam sp_inst_19.INIT_RAM_14 = 256'hF015055FE3555530600055550F0501F50004F020505005105400F143E5500515;
defparam sp_inst_19.INIT_RAM_15 = 256'h505E0F05E0500055F5E3F55E0F0505E50157F300003F005E45351E075F400004;
defparam sp_inst_19.INIT_RAM_16 = 256'hC4200000CCF4C00420C0F4CC00F44F0CF4F04FFF5350055FE35FFF50E5E005E0;
defparam sp_inst_19.INIT_RAM_17 = 256'h3050405220005330C045222000000C4542250000CF4C200CC4FC05330C205330;
defparam sp_inst_19.INIT_RAM_18 = 256'h4FD085020000000F0055000FE35F65402F04FD085020000002F4550042850053;
defparam sp_inst_19.INIT_RAM_19 = 256'h0570F0A0A55460B550750200000705527770010B75771F0C75771F0BF6540CF0;
defparam sp_inst_19.INIT_RAM_1A = 256'hD55FD55500BF350D55460D550750200000705527770010D5FF500F50527153F3;
defparam sp_inst_19.INIT_RAM_1B = 256'h1572577710500205451211101054045EFE40403300FF500F50527153F30570F0;
defparam sp_inst_19.INIT_RAM_1C = 256'h5111055FE3565044FE2FF02750200000057525777104001357F30003F0637121;
defparam sp_inst_19.INIT_RAM_1D = 256'h0055FE35F345C0444552F000005E4505044FEF55F01702005725777104002053;
defparam sp_inst_19.INIT_RAM_1E = 256'hE512F15D5121157257771040020552F4F35251FF354C0555350F02F00D544F15;
defparam sp_inst_19.INIT_RAM_1F = 256'h0F45C0C757710FC40F1E055F5E3F55055FE3F535045EF54504D005454000200F;
defparam sp_inst_19.INIT_RAM_20 = 256'h27F5330571E45C0D5F1C5020057257771030020525F101F45C0DF355B5271121;
defparam sp_inst_19.INIT_RAM_21 = 256'h45C0544F50C050D450CB0D0702000B5275330571F51F2F250A5275330571E555;
defparam sp_inst_19.INIT_RAM_22 = 256'h753305719512110711210C450C951211C545C0100C45C0901211BF35540CB55D;
defparam sp_inst_19.INIT_RAM_23 = 256'h0BFF50DCC5275330571C55B5B45C0B04FEB702000AF354C0801211C45C000B52;
defparam sp_inst_19.INIT_RAM_24 = 256'h000000000049511B000000D705331577F07011005005000FF00043FE85F5D020;
defparam sp_inst_19.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_27 = 256'h400040DBFD020402D1900204E00D520500000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_28 = 256'h40D0410008090859DCE030201304062000960920904304D05040400403E052F6;
defparam sp_inst_19.INIT_RAM_29 = 256'h4040905DF0506D00F346DDC044009346DDC04100C30EDC50C402040D04405020;
defparam sp_inst_19.INIT_RAM_2A = 256'h029D4220C203579D104220C2030309053C20305470540403010B04050C0324F2;
defparam sp_inst_19.INIT_RAM_2B = 256'h0080E9DC00C05002D2007D20550E009D910E0E520F02003FDC0000E410401043;
defparam sp_inst_19.INIT_RAM_2C = 256'h000000000000000000000000000000000000000000000000000000000000050C;
defparam sp_inst_19.INIT_RAM_2D = 256'h0AEF000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2E = 256'h155000880D04455000800AEE115590005D05EA02030004055501139E25A35055;
defparam sp_inst_19.INIT_RAM_2F = 256'h00A80CFA804FA80CF0F30E34D705434D70EC40550EDCC0ED8CC0AC044550AC04;
defparam sp_inst_19.INIT_RAM_30 = 256'h47840784070184010984EF498409CE0403010000700003000000A805D203E001;
defparam sp_inst_19.INIT_RAM_31 = 256'h208700E43D4070F00005009330000958EECF300987095A302490F0C840C0C10F;
defparam sp_inst_19.INIT_RAM_32 = 256'h93F40025FE77035770052E10B240505050633C1F9470ECDC70A3E43D500332C9;
defparam sp_inst_19.INIT_RAM_33 = 256'h4D5A1284A024F5C3024602D050D12547905600640D930D8D940D954A84D340DD;
defparam sp_inst_19.INIT_RAM_34 = 256'h5C9EC108840027E13255084001A104220C255EC770047E204700000000050202;
defparam sp_inst_19.INIT_RAM_35 = 256'h5A89020955A20004277A009191E415505534140403769C6E859C103214891030;
defparam sp_inst_19.INIT_RAM_36 = 256'h0020930EB3020B3A42001DF01550045555A29D4F080202A40255000157004575;
defparam sp_inst_19.INIT_RAM_37 = 256'h8A220E5423D3520EEEE1EEE0EEEE62EEE05C15E5D0EEEEF3EEE0D030AC008502;
defparam sp_inst_19.INIT_RAM_38 = 256'h400000000000000000000000000000000000000000000000000E2E109208A220;
defparam sp_inst_19.INIT_RAM_39 = 256'hE12042E11042E10042E17042E16042E15042E14042E13042E12042E11042E100;
defparam sp_inst_19.INIT_RAM_3A = 256'h5042E14042E13042E12042E11042E10042E17042E16042E15042E14042E13042;
defparam sp_inst_19.INIT_RAM_3B = 256'h42E17042E16042E15042E14042E13042E12042E11042E10042E17042E16042E1;
defparam sp_inst_19.INIT_RAM_3C = 256'h000000000000000000000000000000000000000000000000000000000000022E;
defparam sp_inst_19.INIT_RAM_3D = 256'h0000000000000000000000000000000000005DD0000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_20 (
    .DO({sp_inst_20_dout_w[27:0],sp_inst_20_dout[23:20]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[13],ad[12]}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[23:20]})
);

defparam sp_inst_20.READ_MODE = 1'b0;
defparam sp_inst_20.WRITE_MODE = 2'b01;
defparam sp_inst_20.BIT_WIDTH = 4;
defparam sp_inst_20.BLK_SEL = 3'b010;
defparam sp_inst_20.RESET_MODE = "SYNC";
defparam sp_inst_20.INIT_RAM_00 = 256'h70711111111111180801810190000141417744444477440140184FF801111811;
defparam sp_inst_20.INIT_RAM_01 = 256'h4000110580011777171441BF05980711180840411111111180881011B08800B0;
defparam sp_inst_20.INIT_RAM_02 = 256'hF1090B014F4141441BFF11980711111111111180801810190000117771574417;
defparam sp_inst_20.INIT_RAM_03 = 256'h1001F94144F4414144111109F1090B014F1111111111111180801811090B0101;
defparam sp_inst_20.INIT_RAM_04 = 256'h4F57111F1071111FF141BFF11111F57147401001F58040117177911011777917;
defparam sp_inst_20.INIT_RAM_05 = 256'hF11111B111C111F41174F1904F111111111111180801810190014F4174F14174;
defparam sp_inst_20.INIT_RAM_06 = 256'h5714174F11F41740F141174F8F8711114F111111C111F1090B014F111111C111;
defparam sp_inst_20.INIT_RAM_07 = 256'h111C111F4174F41174F11111071111F111114FBB10004F4174F141744F81111F;
defparam sp_inst_20.INIT_RAM_08 = 256'h111F5711F1F410741F41174F41744F81BFF71111F574174F811111F41074F111;
defparam sp_inst_20.INIT_RAM_09 = 256'h14409047711B411044090477444F191F4174141B1F1111F4174141B1F111111C;
defparam sp_inst_20.INIT_RAM_0A = 256'hF5714F119991BF074040180808F8111101177711191F8180A10808001814110B;
defparam sp_inst_20.INIT_RAM_0B = 256'h9811F8184F8981014F111B011888B00B001F18111B088800B001401171771111;
defparam sp_inst_20.INIT_RAM_0C = 256'h0211B00B10414412022026414411B1008BF9BB10011777191710F8184F8181F8;
defparam sp_inst_20.INIT_RAM_0D = 256'h00B10144202120208111100141411111164111101616441441B00B1014620212;
defparam sp_inst_20.INIT_RAM_0E = 256'h19991BF07404081000B10111110146411411111146141B00B10146202120211B;
defparam sp_inst_20.INIT_RAM_0F = 256'h4111111B1C119F8F81F11474F118711180840141111119084081187771571401;
defparam sp_inst_20.INIT_RAM_10 = 256'h4F1F148C7F84F1FF4FFF4F41444F4F1000B1111FF11111B8F11111B84FF184F1;
defparam sp_inst_20.INIT_RAM_11 = 256'h401411111198BBF14FFF11B114F14F1F11108180BF814F14C87F84F1B1114FF1;
defparam sp_inst_20.INIT_RAM_12 = 256'h00101041000414177797FF184F14111111B1C119F8FFF1FF11474F1187111808;
defparam sp_inst_20.INIT_RAM_13 = 256'h4409047744FF1FF114BF11BF100F4F114B0FF1F0111B401801114B0041001001;
defparam sp_inst_20.INIT_RAM_14 = 256'hB001011777111108080811114F818091408090081814110B14409047711B4101;
defparam sp_inst_20.INIT_RAM_15 = 256'h181F8981F81840117177911F898101F1B111B088800B001F417117B11B088800;
defparam sp_inst_20.INIT_RAM_16 = 256'h1411141111641144111164118064468164684BF9171001177719BB10F1F881F8;
defparam sp_inst_20.INIT_RAM_17 = 256'h1114411111111111114111111141114141114114164111111461111111111111;
defparam sp_inst_20.INIT_RAM_18 = 256'h1BF071118084040808118887771571440991BF07111808404084114440714111;
defparam sp_inst_20.INIT_RAM_19 = 256'hC119F8F8F11474F118711180840141111119018F11111B8F11111B8F57144F99;
defparam sp_inst_20.INIT_RAM_1A = 256'hF119F11108F9710F11474F118711180840141111119018F1FF184F14111111B1;
defparam sp_inst_20.INIT_RAM_1B = 256'h11111111180801810100001C041444179744447744FF184F14111111B1C119F8;
defparam sp_inst_20.INIT_RAM_1C = 256'h1000011777171441BF05980711180840411111111180881011B08800B0707111;
defparam sp_inst_20.INIT_RAM_1D = 256'h4011777157417400011058000A1F4141441BFF11980711111111111180801810;
defparam sp_inst_20.INIT_RAM_1E = 256'hF100B01F111111111111180801811090B01011F571474010010580FC4F100B01;
defparam sp_inst_20.INIT_RAM_1F = 256'h4F4174F111114FF14B1F01171779110117779171001F914144F4414144111109;
defparam sp_inst_20.INIT_RAM_20 = 256'h11B111C111F4174F190F11111111111118080181019001F4174F5711F1071111;
defparam sp_inst_20.INIT_RAM_21 = 256'h4174141B107410F4147F8F8711114F111111C111F1090B014F111111C111F111;
defparam sp_inst_20.INIT_RAM_22 = 256'h1111C111F111110711114F4147F11111F14174004F4174F81111F5711447F11F;
defparam sp_inst_20.INIT_RAM_23 = 256'h1FBB10F7F111111C111F11F1F4174F81BFF711114F571474F81111F417044F11;
defparam sp_inst_20.INIT_RAM_24 = 256'h0000000000633326000008AC01111111A01811991001401BF0904787F191F111;
defparam sp_inst_20.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_27 = 256'h6203602662032723346203366200272620000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_28 = 256'h6062630007060767266030306503054033033033007404405040603606602757;
defparam sp_inst_20.INIT_RAM_29 = 256'h7072606560707500676665626300776665626300660363606627260626306272;
defparam sp_inst_20.INIT_RAM_2A = 256'h0765677733066765626777330606760673306066606707077606072606077767;
defparam sp_inst_20.INIT_RAM_2B = 256'h0070665670606707577075776606706566060666060770753670703760706066;
defparam sp_inst_20.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000504;
defparam sp_inst_20.INIT_RAM_2D = 256'h0066000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2E = 256'h3670307706263670303300636367500026026027040206266702666654072022;
defparam sp_inst_20.INIT_RAM_2F = 256'h2207265072550726506706766506776650336267026660267660062636700626;
defparam sp_inst_20.INIT_RAM_30 = 256'h6767076507066506066525666706660307032223322233222322072233076224;
defparam sp_inst_20.INIT_RAM_31 = 256'h7266202776727262227722066222206636366220672673707740606650606625;
defparam sp_inst_20.INIT_RAM_32 = 256'h7767007766670777620272676750202020777236766233666206277662077736;
defparam sp_inst_20.INIT_RAM_33 = 256'h6220676702376667076707676006767662667267006726626700667366277006;
defparam sp_inst_20.INIT_RAM_34 = 256'h6363340777207636636707603606267773367337620662727700000000023303;
defparam sp_inst_20.INIT_RAM_35 = 256'h7076032667077007767052434437667067633626063622722522324334244270;
defparam sp_inst_20.INIT_RAM_36 = 256'h7072660666072660677066606660266667076366260727062767000667026676;
defparam sp_inst_20.INIT_RAM_37 = 256'h7377027776676702222422202222442220266667202222552220026236207227;
defparam sp_inst_20.INIT_RAM_38 = 256'h7000000000000000000000000000000000000000000000000002766267073770;
defparam sp_inst_20.INIT_RAM_39 = 256'h6737776737776737776737776737776737776737776737776737776737776737;
defparam sp_inst_20.INIT_RAM_3A = 256'h3777673777673777673777673777673777673777673777673777673777673777;
defparam sp_inst_20.INIT_RAM_3B = 256'h7767377767377767377767377767377767377767377767377767377767377767;
defparam sp_inst_20.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000776;
defparam sp_inst_20.INIT_RAM_3D = 256'h00000000000000000000000000000000000006C0000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_21 (
    .DO({sp_inst_21_dout_w[27:0],sp_inst_21_dout[27:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[13],ad[12]}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[27:24]})
);

defparam sp_inst_21.READ_MODE = 1'b0;
defparam sp_inst_21.WRITE_MODE = 2'b01;
defparam sp_inst_21.BIT_WIDTH = 4;
defparam sp_inst_21.BLK_SEL = 3'b010;
defparam sp_inst_21.RESET_MODE = "SYNC";
defparam sp_inst_21.INIT_RAM_00 = 256'h0000000000000002020020802404800000000000000033C03C023372C0000200;
defparam sp_inst_21.INIT_RAM_01 = 256'h0404004324C00000000000358322000002823030000000002022000024220420;
defparam sp_inst_21.INIT_RAM_02 = 256'h3082020033000030035B0022000000000000002020020802404C000000303000;
defparam sp_inst_21.INIT_RAM_03 = 256'h0400F20000733000000000823082020033000000000000002020020082020040;
defparam sp_inst_21.INIT_RAM_04 = 256'h333000070400000370303570000033000004004073243C000000200C00000200;
defparam sp_inst_21.INIT_RAM_05 = 256'h30000020003000300000F0243300000000000002020020802400330000300000;
defparam sp_inst_21.INIT_RAM_06 = 256'h3000000300300004300000032320000033000000300030820200330000003000;
defparam sp_inst_21.INIT_RAM_07 = 256'h0003000300003000003000000000003000003323044433000030000033200003;
defparam sp_inst_21.INIT_RAM_08 = 256'h0003300070300400030000030000332035300000330000032000003004003000;
defparam sp_inst_21.INIT_RAM_09 = 256'h0008200000020004008200003333020300000002030000300000002030000003;
defparam sp_inst_21.INIT_RAM_0A = 256'h33000300222035000434028282B20000C00000000203203420C802C802000042;
defparam sp_inst_21.INIT_RAM_0B = 256'h22003203332220403300024002222042000302000242220420003C0000000000;
defparam sp_inst_21.INIT_RAM_0C = 256'hC0002C820C000000C00C00000000208892322304C00000020004320333202032;
defparam sp_inst_21.INIT_RAM_0D = 256'hC820C0000C000C0820000880000000000000000400000000302C820C0000C000;
defparam sp_inst_21.INIT_RAM_0E = 256'h02220350004343088820C0000040000000000000000002C820C0000C000C0002;
defparam sp_inst_21.INIT_RAM_0F = 256'h3000000203002723203000007002000028230030000002423C20080000300000;
defparam sp_inst_21.INIT_RAM_10 = 256'h330300232B2330FF333F3300000B33088C20000F300000223000002233F02330;
defparam sp_inst_21.INIT_RAM_11 = 256'h300300000022223033FF0020003033030004202023203300322B233020003F30;
defparam sp_inst_21.INIT_RAM_12 = 256'h000404204880000000203F023303000000203002723730B30000070020000282;
defparam sp_inst_21.INIT_RAM_13 = 256'h00820000333F0B300223002F088333002243707C00023C02C000228420440C40;
defparam sp_inst_21.INIT_RAM_14 = 256'h2000C000000000C282820000332034203C802C82020000420008200000020040;
defparam sp_inst_21.INIT_RAM_15 = 256'h0203222032033C00000020032220403020002422204200070000002002422204;
defparam sp_inst_21.INIT_RAM_16 = 256'h00000000000000000000000094000090000902320004C0000002230430323032;
defparam sp_inst_21.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_18 = 256'h0350000028230342C20088800003000002203500000282303420000300000000;
defparam sp_inst_21.INIT_RAM_19 = 256'h3002723230000070020000282300300000024023000002230000022330000322;
defparam sp_inst_21.INIT_RAM_1A = 256'h3002300042320043000007002000028230030000002402303F02330300000020;
defparam sp_inst_21.INIT_RAM_1B = 256'h0000000002020020804048038000000020000000333F02330300000020300272;
defparam sp_inst_21.INIT_RAM_1C = 256'h0404C00000000000358322000002823030000000002022000024220420000000;
defparam sp_inst_21.INIT_RAM_1D = 256'h3C00000030000040400432480203000030035B00220000000000000020200208;
defparam sp_inst_21.INIT_RAM_1E = 256'h308020030000000000000202002008202004003300000400404324F333080200;
defparam sp_inst_21.INIT_RAM_1F = 256'h33000030000033703305C000000200C000002000400F20000073300000000082;
defparam sp_inst_21.INIT_RAM_20 = 256'h002000300030000F024300000000000002020020802400300003300070400000;
defparam sp_inst_21.INIT_RAM_21 = 256'h0000000200000030000323200000330000003000308202003300000030003000;
defparam sp_inst_21.INIT_RAM_22 = 256'h0000300030000000000033000030000030000004330000320000330000003003;
defparam sp_inst_21.INIT_RAM_23 = 256'h0323043030000003000300703000032035300000333000003200003000403300;
defparam sp_inst_21.INIT_RAM_24 = 256'hCCCCCCCCC05162A50000C88CC00000002002002204C03C034424002030203000;
defparam sp_inst_21.INIT_RAM_25 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam sp_inst_21.INIT_RAM_26 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam sp_inst_21.INIT_RAM_27 = 256'h020840DD0D08014804340884340A00192CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam sp_inst_21.INIT_RAM_28 = 256'h50EC4000090405A4D0404040C504011099095091000F0F5000F000840BF02D19;
defparam sp_inst_21.INIT_RAM_29 = 256'h90D4D040503010002349F05C40004349F05C40009D0D13C00075150EC4000251;
defparam sp_inst_21.INIT_RAM_2A = 256'h052045E1330202204C45E1330701220E30300037003305040B050D4C01040920;
defparam sp_inst_21.INIT_RAM_2B = 256'h00404F019010190409902019020990E0E2090E4100019086E19090D040404030;
defparam sp_inst_21.INIT_RAM_2C = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC0C0C;
defparam sp_inst_21.INIT_RAM_2D = 256'h0A4DCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam sp_inst_21.INIT_RAM_2E = 256'h0A3080A50EC40A3020880D5040A300004004005004000ECCA301EFE4A2093032;
defparam sp_inst_21.INIT_RAM_2F = 256'h3005D4005D8F05D0302504401D041401D0AE2CA30E2050E20050D5C40A30D5C4;
defparam sp_inst_21.INIT_RAM_30 = 256'hFE0F0E0F0E0E0F0E040F04F40F040404060A00080000400000000508040A4004;
defparam sp_inst_21.INIT_RAM_31 = 256'h9C0550AE4508035009F30091840A00C10F47840AEECE3010F0E070C0F0C0EEC4;
defparam sp_inst_21.INIT_RAM_32 = 256'h0005001D6702050155047E2050904040401EC2A405550351550A1E450305E433;
defparam sp_inst_21.INIT_RAM_33 = 256'hD5007005087F304801010D5130AC54F5E9E25A050AE54A84050AD4F3A4D050A5;
defparam sp_inst_21.INIT_RAM_34 = 256'h3460340D5120E1C483A305208404C45E133A3034550A3E4354CCCC0000002404;
defparam sp_inst_21.INIT_RAM_35 = 256'h30540ECEA3029005102092F004004A305C10A209019C60205460E819C3104850;
defparam sp_inst_21.INIT_RAM_36 = 256'h90432F0508043F80F12020702020A402A30D151255043502C5A30002020A402A;
defparam sp_inst_21.INIT_RAM_37 = 256'hA0540A050C50290AEEE4EEE0EEEE11EEE08AE943D0EEEE9FEEE0A0A609C0A852;
defparam sp_inst_21.INIT_RAM_38 = 256'h9CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC0E5423D50A0540;
defparam sp_inst_21.INIT_RAM_39 = 256'h4FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9;
defparam sp_inst_21.INIT_RAM_3A = 256'hF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF990;
defparam sp_inst_21.INIT_RAM_3B = 256'hF04FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904FF9904F;
defparam sp_inst_21.INIT_RAM_3C = 256'h00000C0000000000000000C00C00CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC0404;
defparam sp_inst_21.INIT_RAM_3D = 256'h00000000000000000000000000000000000006B0000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_22 (
    .DO({sp_inst_22_dout_w[27:0],sp_inst_22_dout[31:28]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[13],ad[12]}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:28]})
);

defparam sp_inst_22.READ_MODE = 1'b0;
defparam sp_inst_22.WRITE_MODE = 2'b01;
defparam sp_inst_22.BIT_WIDTH = 4;
defparam sp_inst_22.BLK_SEL = 3'b010;
defparam sp_inst_22.RESET_MODE = "SYNC";
defparam sp_inst_22.INIT_RAM_00 = 256'h0400000000000000606000500146500000000000000000400400054040000000;
defparam sp_inst_22.INIT_RAM_01 = 256'h0444004004400000000000015000400000500400000000000600060006000400;
defparam sp_inst_22.INIT_RAM_02 = 256'h5050404005000000001500004000000000000006060005001464000000000000;
defparam sp_inst_22.INIT_RAM_03 = 256'h0140500000400000000000505050404005000000000000000606000050404040;
defparam sp_inst_22.INIT_RAM_04 = 256'h0500000404000005400001600000500000040440400404000000000400000000;
defparam sp_inst_22.INIT_RAM_05 = 256'h5000000000000050000050010500000000000000606000500140050000500000;
defparam sp_inst_22.INIT_RAM_06 = 256'h0000000400500004500000050400000005000000000050504040050000000000;
defparam sp_inst_22.INIT_RAM_07 = 256'h0000000500005000005000004000005000000500014405000050000005000005;
defparam sp_inst_22.INIT_RAM_08 = 256'h0005000040500400050000050000050001400000500000050000005004005000;
defparam sp_inst_22.INIT_RAM_09 = 256'h0005040000000001005040000005000500000000050000500000000050000000;
defparam sp_inst_22.INIT_RAM_0A = 256'h5000060000000140040600505050000040000000000500040042001600000010;
defparam sp_inst_22.INIT_RAM_0B = 256'h0000500005000040050000600000004004050000006000040040040000000000;
defparam sp_inst_22.INIT_RAM_0C = 256'h5000066006000000500500000000005620500001400000000001500005000050;
defparam sp_inst_22.INIT_RAM_0D = 256'h6600600005000505000005600000000000000001000000000006600600005000;
defparam sp_inst_22.INIT_RAM_0E = 256'h0000001400406005660060000010000000000000000000660060000500050000;
defparam sp_inst_22.INIT_RAM_0F = 256'h0000000000000606005000004000000005004000000000400400020000000060;
defparam sp_inst_22.INIT_RAM_10 = 256'h0505000005005065054505000006050566000006500000005000000005500040;
defparam sp_inst_22.INIT_RAM_11 = 256'h0400000000000050055500000050050500060004060005000005005000000650;
defparam sp_inst_22.INIT_RAM_12 = 256'h5404040045500000000055000400000000000000605450650000040000000050;
defparam sp_inst_22.INIT_RAM_13 = 256'h0050400000560650000500060566050000654044000004004000005400440540;
defparam sp_inst_22.INIT_RAM_14 = 256'h0040400000000050505000000500040004200160000000100005040000000010;
defparam sp_inst_22.INIT_RAM_15 = 256'h0005000050000400000000050000405000000600004004040000000000600004;
defparam sp_inst_22.INIT_RAM_16 = 256'h0000000000000000000000002100002000020050000140000000000150500050;
defparam sp_inst_22.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_18 = 256'h0014000005004060400022200000000060000140000050040600000004000000;
defparam sp_inst_22.INIT_RAM_19 = 256'h0000606050000040000000050040000000004005000000050000000500000600;
defparam sp_inst_22.INIT_RAM_1A = 256'h5000500060500015000004000000005004000000000400505500040000000000;
defparam sp_inst_22.INIT_RAM_1B = 256'h0000000000606000501465005000000000000000005500040000000000000060;
defparam sp_inst_22.INIT_RAM_1C = 256'h0146400000000000015000400000500400000000000600060006000400040000;
defparam sp_inst_22.INIT_RAM_1D = 256'h0400000000000044400400454005000000001500004000000000000006060005;
defparam sp_inst_22.INIT_RAM_1E = 256'h5054040500000000000000606000050404040050000004044040045005054040;
defparam sp_inst_22.INIT_RAM_1F = 256'h0500005000000540000140000000004000000000140500000040000000000050;
defparam sp_inst_22.INIT_RAM_20 = 256'h0000000000500005001500000000000000606000500140500005000040400000;
defparam sp_inst_22.INIT_RAM_21 = 256'h0000000004000450000504000000050000000000505040400500000000005000;
defparam sp_inst_22.INIT_RAM_22 = 256'h0000000050000040000005000050000050000044050000500000500000004005;
defparam sp_inst_22.INIT_RAM_23 = 256'h0500015050000000000500405000050001400000050000005000005000400500;
defparam sp_inst_22.INIT_RAM_24 = 256'h1111111110663306000042214000000006000000014004001606000050005000;
defparam sp_inst_22.INIT_RAM_25 = 256'h1111111111111111111111111111111111111111111111111111111111111111;
defparam sp_inst_22.INIT_RAM_26 = 256'h1111111111111111111111111111111111111111111111111111111111111111;
defparam sp_inst_22.INIT_RAM_27 = 256'h2707602222073657366407767700326671111111111111111111111111111111;
defparam sp_inst_22.INIT_RAM_28 = 256'h7033620006070235207060606706066003303303302606705060007606603346;
defparam sp_inst_22.INIT_RAM_29 = 256'h6057607070603000776760736200776760736200660566607076670336200666;
defparam sp_inst_22.INIT_RAM_2A = 256'h0630663666070730736636660706730367607076007606072606057606072670;
defparam sp_inst_22.INIT_RAM_2B = 256'h0070760660606606066070660706606067060376070670663660705270606060;
defparam sp_inst_22.INIT_RAM_2C = 256'h1111111111111111111111111111111111111111111111111111111111110404;
defparam sp_inst_22.INIT_RAM_2D = 256'h0066111111111111111111111111111111111111111111111111111111111111;
defparam sp_inst_22.INIT_RAM_2E = 256'h2370303203362370307700726237400062062023040003363702666635007073;
defparam sp_inst_22.INIT_RAM_2F = 256'h4202355023640232407606726406672640067337026260262260073623700736;
defparam sp_inst_22.INIT_RAM_30 = 256'h6626062606062606072607672607070607002233222332223322022326007227;
defparam sp_inst_22.INIT_RAM_31 = 256'h6376500276260772206622066720226625676720363662606260706260603637;
defparam sp_inst_22.INIT_RAM_32 = 256'h2726002666270676650662726260606060632336266507666503627626063776;
defparam sp_inst_22.INIT_RAM_33 = 256'h2230622604367266062600666006676666677326006673662600676736626006;
defparam sp_inst_22.INIT_RAM_34 = 256'h7772740026703636663702707707366366637076650062776611110000033606;
defparam sp_inst_22.INIT_RAM_35 = 256'h7026033637077006627043423422737026603336062272733552224224334260;
defparam sp_inst_22.INIT_RAM_36 = 256'h7077760626077660667072607270062737036267660776073637000727006273;
defparam sp_inst_22.INIT_RAM_37 = 256'h0367007626627600222422202222442220736776202222442220023626300727;
defparam sp_inst_22.INIT_RAM_38 = 256'h6111111111111111111111111111111111111111111111111102777666003670;
defparam sp_inst_22.INIT_RAM_39 = 256'h6556606556606556606556606556606556606556606556606556606556606556;
defparam sp_inst_22.INIT_RAM_3A = 256'h5660655660655660655660655660655660655660655660655660655660655660;
defparam sp_inst_22.INIT_RAM_3B = 256'h5065566065566065566065566065566065566065566065566065566065566065;
defparam sp_inst_22.INIT_RAM_3C = 256'h0000010000000008880080188100111111111111111111111111111111110706;
defparam sp_inst_22.INIT_RAM_3D = 256'h0000000000000000000000000000000000000EA0000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_23 (
    .DO(sp_inst_23_dout[31:0]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[8:0],gw_gnd,gw_vcc,gw_vcc,gw_vcc,gw_vcc}),
    .DI(din[31:0])
);

defparam sp_inst_23.READ_MODE = 1'b0;
defparam sp_inst_23.WRITE_MODE = 2'b01;
defparam sp_inst_23.BIT_WIDTH = 32;
defparam sp_inst_23.BLK_SEL = 3'b001;
defparam sp_inst_23.RESET_MODE = "SYNC";
defparam sp_inst_23.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(spx9_inst_0_dout[0]),
  .I1(spx9_inst_1_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(spx9_inst_2_dout[0]),
  .I1(spx9_inst_3_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_1)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(sp_inst_15_dout[0]),
  .I1(sp_inst_23_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_18 (
  .O(dout[0]),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_0)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(spx9_inst_0_dout[1]),
  .I1(spx9_inst_1_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(spx9_inst_2_dout[1]),
  .I1(spx9_inst_3_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(mux_o_31),
  .I1(mux_o_32),
  .S0(dff_q_1)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(sp_inst_15_dout[1]),
  .I1(sp_inst_23_dout[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_37 (
  .O(dout[1]),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_0)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(spx9_inst_0_dout[2]),
  .I1(spx9_inst_1_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(spx9_inst_2_dout[2]),
  .I1(spx9_inst_3_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_50),
  .I1(mux_o_51),
  .S0(dff_q_1)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(sp_inst_15_dout[2]),
  .I1(sp_inst_23_dout[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_56 (
  .O(dout[2]),
  .I0(mux_o_54),
  .I1(mux_o_55),
  .S0(dff_q_0)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(spx9_inst_0_dout[3]),
  .I1(spx9_inst_1_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(spx9_inst_2_dout[3]),
  .I1(spx9_inst_3_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_69),
  .I1(mux_o_70),
  .S0(dff_q_1)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(sp_inst_15_dout[3]),
  .I1(sp_inst_23_dout[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_75 (
  .O(dout[3]),
  .I0(mux_o_73),
  .I1(mux_o_74),
  .S0(dff_q_0)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(spx9_inst_0_dout[4]),
  .I1(spx9_inst_1_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(spx9_inst_2_dout[4]),
  .I1(spx9_inst_3_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(dff_q_1)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(sp_inst_16_dout[4]),
  .I1(sp_inst_23_dout[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_94 (
  .O(dout[4]),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(dff_q_0)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(spx9_inst_0_dout[5]),
  .I1(spx9_inst_1_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(spx9_inst_2_dout[5]),
  .I1(spx9_inst_3_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_1)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(sp_inst_16_dout[5]),
  .I1(sp_inst_23_dout[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_113 (
  .O(dout[5]),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(dff_q_0)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(spx9_inst_0_dout[6]),
  .I1(spx9_inst_1_dout[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(spx9_inst_2_dout[6]),
  .I1(spx9_inst_3_dout[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_1)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(sp_inst_16_dout[6]),
  .I1(sp_inst_23_dout[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_132 (
  .O(dout[6]),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_0)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(spx9_inst_0_dout[7]),
  .I1(spx9_inst_1_dout[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(spx9_inst_2_dout[7]),
  .I1(spx9_inst_3_dout[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_145),
  .I1(mux_o_146),
  .S0(dff_q_1)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(sp_inst_16_dout[7]),
  .I1(sp_inst_23_dout[7]),
  .S0(dff_q_1)
);
MUX2 mux_inst_151 (
  .O(dout[7]),
  .I0(mux_o_149),
  .I1(mux_o_150),
  .S0(dff_q_0)
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(spx9_inst_0_dout[8]),
  .I1(spx9_inst_1_dout[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(spx9_inst_2_dout[8]),
  .I1(spx9_inst_3_dout[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(mux_o_164),
  .I1(mux_o_165),
  .S0(dff_q_1)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(sp_inst_17_dout[8]),
  .I1(sp_inst_23_dout[8]),
  .S0(dff_q_1)
);
MUX2 mux_inst_170 (
  .O(dout[8]),
  .I0(mux_o_168),
  .I1(mux_o_169),
  .S0(dff_q_0)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(spx9_inst_4_dout[9]),
  .I1(spx9_inst_5_dout[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(spx9_inst_6_dout[9]),
  .I1(spx9_inst_7_dout[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(dff_q_1)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(sp_inst_17_dout[9]),
  .I1(sp_inst_23_dout[9]),
  .S0(dff_q_1)
);
MUX2 mux_inst_189 (
  .O(dout[9]),
  .I0(mux_o_187),
  .I1(mux_o_188),
  .S0(dff_q_0)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(spx9_inst_4_dout[10]),
  .I1(spx9_inst_5_dout[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(spx9_inst_6_dout[10]),
  .I1(spx9_inst_7_dout[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_202),
  .I1(mux_o_203),
  .S0(dff_q_1)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(sp_inst_17_dout[10]),
  .I1(sp_inst_23_dout[10]),
  .S0(dff_q_1)
);
MUX2 mux_inst_208 (
  .O(dout[10]),
  .I0(mux_o_206),
  .I1(mux_o_207),
  .S0(dff_q_0)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(spx9_inst_4_dout[11]),
  .I1(spx9_inst_5_dout[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(spx9_inst_6_dout[11]),
  .I1(spx9_inst_7_dout[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_1)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(sp_inst_17_dout[11]),
  .I1(sp_inst_23_dout[11]),
  .S0(dff_q_1)
);
MUX2 mux_inst_227 (
  .O(dout[11]),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(dff_q_0)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(spx9_inst_4_dout[12]),
  .I1(spx9_inst_5_dout[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(spx9_inst_6_dout[12]),
  .I1(spx9_inst_7_dout[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_240),
  .I1(mux_o_241),
  .S0(dff_q_1)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(sp_inst_18_dout[12]),
  .I1(sp_inst_23_dout[12]),
  .S0(dff_q_1)
);
MUX2 mux_inst_246 (
  .O(dout[12]),
  .I0(mux_o_244),
  .I1(mux_o_245),
  .S0(dff_q_0)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(spx9_inst_4_dout[13]),
  .I1(spx9_inst_5_dout[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(spx9_inst_6_dout[13]),
  .I1(spx9_inst_7_dout[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(mux_o_259),
  .I1(mux_o_260),
  .S0(dff_q_1)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(sp_inst_18_dout[13]),
  .I1(sp_inst_23_dout[13]),
  .S0(dff_q_1)
);
MUX2 mux_inst_265 (
  .O(dout[13]),
  .I0(mux_o_263),
  .I1(mux_o_264),
  .S0(dff_q_0)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(spx9_inst_4_dout[14]),
  .I1(spx9_inst_5_dout[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(spx9_inst_6_dout[14]),
  .I1(spx9_inst_7_dout[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(dff_q_1)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(sp_inst_18_dout[14]),
  .I1(sp_inst_23_dout[14]),
  .S0(dff_q_1)
);
MUX2 mux_inst_284 (
  .O(dout[14]),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_0)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(spx9_inst_4_dout[15]),
  .I1(spx9_inst_5_dout[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(spx9_inst_6_dout[15]),
  .I1(spx9_inst_7_dout[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_297),
  .I1(mux_o_298),
  .S0(dff_q_1)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(sp_inst_18_dout[15]),
  .I1(sp_inst_23_dout[15]),
  .S0(dff_q_1)
);
MUX2 mux_inst_303 (
  .O(dout[15]),
  .I0(mux_o_301),
  .I1(mux_o_302),
  .S0(dff_q_0)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(spx9_inst_4_dout[16]),
  .I1(spx9_inst_5_dout[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(spx9_inst_6_dout[16]),
  .I1(spx9_inst_7_dout[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(mux_o_316),
  .I1(mux_o_317),
  .S0(dff_q_1)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(sp_inst_19_dout[16]),
  .I1(sp_inst_23_dout[16]),
  .S0(dff_q_1)
);
MUX2 mux_inst_322 (
  .O(dout[16]),
  .I0(mux_o_320),
  .I1(mux_o_321),
  .S0(dff_q_0)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(spx9_inst_4_dout[17]),
  .I1(spx9_inst_5_dout[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(spx9_inst_6_dout[17]),
  .I1(spx9_inst_7_dout[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_335),
  .I1(mux_o_336),
  .S0(dff_q_1)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(sp_inst_19_dout[17]),
  .I1(sp_inst_23_dout[17]),
  .S0(dff_q_1)
);
MUX2 mux_inst_341 (
  .O(dout[17]),
  .I0(mux_o_339),
  .I1(mux_o_340),
  .S0(dff_q_0)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(sp_inst_19_dout[18]),
  .I1(sp_inst_23_dout[18]),
  .S0(dff_q_1)
);
MUX2 mux_inst_353 (
  .O(dout[18]),
  .I0(sp_inst_8_dout[18]),
  .I1(mux_o_352),
  .S0(dff_q_0)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(sp_inst_19_dout[19]),
  .I1(sp_inst_23_dout[19]),
  .S0(dff_q_1)
);
MUX2 mux_inst_365 (
  .O(dout[19]),
  .I0(sp_inst_8_dout[19]),
  .I1(mux_o_364),
  .S0(dff_q_0)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(sp_inst_20_dout[20]),
  .I1(sp_inst_23_dout[20]),
  .S0(dff_q_1)
);
MUX2 mux_inst_377 (
  .O(dout[20]),
  .I0(sp_inst_9_dout[20]),
  .I1(mux_o_376),
  .S0(dff_q_0)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(sp_inst_20_dout[21]),
  .I1(sp_inst_23_dout[21]),
  .S0(dff_q_1)
);
MUX2 mux_inst_389 (
  .O(dout[21]),
  .I0(sp_inst_9_dout[21]),
  .I1(mux_o_388),
  .S0(dff_q_0)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(sp_inst_20_dout[22]),
  .I1(sp_inst_23_dout[22]),
  .S0(dff_q_1)
);
MUX2 mux_inst_401 (
  .O(dout[22]),
  .I0(sp_inst_10_dout[22]),
  .I1(mux_o_400),
  .S0(dff_q_0)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(sp_inst_20_dout[23]),
  .I1(sp_inst_23_dout[23]),
  .S0(dff_q_1)
);
MUX2 mux_inst_413 (
  .O(dout[23]),
  .I0(sp_inst_10_dout[23]),
  .I1(mux_o_412),
  .S0(dff_q_0)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(sp_inst_21_dout[24]),
  .I1(sp_inst_23_dout[24]),
  .S0(dff_q_1)
);
MUX2 mux_inst_425 (
  .O(dout[24]),
  .I0(sp_inst_11_dout[24]),
  .I1(mux_o_424),
  .S0(dff_q_0)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(sp_inst_21_dout[25]),
  .I1(sp_inst_23_dout[25]),
  .S0(dff_q_1)
);
MUX2 mux_inst_437 (
  .O(dout[25]),
  .I0(sp_inst_11_dout[25]),
  .I1(mux_o_436),
  .S0(dff_q_0)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(sp_inst_21_dout[26]),
  .I1(sp_inst_23_dout[26]),
  .S0(dff_q_1)
);
MUX2 mux_inst_449 (
  .O(dout[26]),
  .I0(sp_inst_12_dout[26]),
  .I1(mux_o_448),
  .S0(dff_q_0)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(sp_inst_21_dout[27]),
  .I1(sp_inst_23_dout[27]),
  .S0(dff_q_1)
);
MUX2 mux_inst_461 (
  .O(dout[27]),
  .I0(sp_inst_12_dout[27]),
  .I1(mux_o_460),
  .S0(dff_q_0)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(sp_inst_22_dout[28]),
  .I1(sp_inst_23_dout[28]),
  .S0(dff_q_1)
);
MUX2 mux_inst_473 (
  .O(dout[28]),
  .I0(sp_inst_13_dout[28]),
  .I1(mux_o_472),
  .S0(dff_q_0)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(sp_inst_22_dout[29]),
  .I1(sp_inst_23_dout[29]),
  .S0(dff_q_1)
);
MUX2 mux_inst_485 (
  .O(dout[29]),
  .I0(sp_inst_13_dout[29]),
  .I1(mux_o_484),
  .S0(dff_q_0)
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(sp_inst_22_dout[30]),
  .I1(sp_inst_23_dout[30]),
  .S0(dff_q_1)
);
MUX2 mux_inst_497 (
  .O(dout[30]),
  .I0(sp_inst_14_dout[30]),
  .I1(mux_o_496),
  .S0(dff_q_0)
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(sp_inst_22_dout[31]),
  .I1(sp_inst_23_dout[31]),
  .S0(dff_q_1)
);
MUX2 mux_inst_509 (
  .O(dout[31]),
  .I0(sp_inst_14_dout[31]),
  .I1(mux_o_508),
  .S0(dff_q_0)
);
endmodule //Gowin_SP_Instr
